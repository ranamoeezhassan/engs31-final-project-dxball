library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity game_win_rom is
  Port (
    clk        : in  std_logic;
    row        : in  std_logic_vector(7 downto 0);
    col        : in  std_logic_vector(6 downto 0);
    color_data : out std_logic_vector(11 downto 0)
  );
end entity;

architecture Behavioral of game_win_rom is
  signal addr : std_logic_vector(14 downto 0);
  signal row_reg : std_logic_vector(7 downto 0);
  signal  col_reg : std_logic_vector(6 downto 0);
begin

  process(clk)
  begin
    if rising_edge(clk) then
      row_reg <= row;
      col_reg <= col;
    end if;
  end process;

  addr <= row_reg & col_reg;

  process(addr)
  begin
    case addr is
      when "000000000000000" => color_data <= "000000000000";
      when "000000000000001" => color_data <= "000000000000";
      when "000000000000010" => color_data <= "000000000000";
      when "000000000000011" => color_data <= "000000000000";
      when "000000000000100" => color_data <= "000000000000";
      when "000000000000101" => color_data <= "000000000000";
      when "000000000000110" => color_data <= "000000000000";
      when "000000000000111" => color_data <= "000000000000";
      when "000000000001000" => color_data <= "000000000000";
      when "000000000001001" => color_data <= "000000000000";
      when "000000000001010" => color_data <= "000000000000";
      when "000000000001011" => color_data <= "000000000000";
      when "000000000001100" => color_data <= "000000000000";
      when "000000000001101" => color_data <= "000000000000";
      when "000000000001110" => color_data <= "000000000000";
      when "000000000001111" => color_data <= "000000000000";
      when "000000000010000" => color_data <= "000000000000";
      when "000000000010001" => color_data <= "000000000000";
      when "000000000010010" => color_data <= "000000000000";
      when "000000000010011" => color_data <= "000000000000";
      when "000000000010100" => color_data <= "000000000000";
      when "000000000010101" => color_data <= "000000000000";
      when "000000000010110" => color_data <= "000000000000";
      when "000000000010111" => color_data <= "000000000000";
      when "000000000011000" => color_data <= "000000000000";
      when "000000000011001" => color_data <= "000000000000";
      when "000000000011010" => color_data <= "000000000000";
      when "000000000011011" => color_data <= "000000000000";
      when "000000000011100" => color_data <= "000000000000";
      when "000000000011101" => color_data <= "000000000000";
      when "000000000011110" => color_data <= "000000000000";
      when "000000000011111" => color_data <= "000000000000";
      when "000000000100000" => color_data <= "000000000000";
      when "000000000100001" => color_data <= "000000000000";
      when "000000000100010" => color_data <= "000000000000";
      when "000000000100011" => color_data <= "000000000000";
      when "000000000100100" => color_data <= "000000000000";
      when "000000000100101" => color_data <= "000000000000";
      when "000000000100110" => color_data <= "000000000000";
      when "000000000100111" => color_data <= "000000000000";
      when "000000000101000" => color_data <= "000000000000";
      when "000000000101001" => color_data <= "000000000000";
      when "000000000101010" => color_data <= "000000000000";
      when "000000000101011" => color_data <= "000000000000";
      when "000000000101100" => color_data <= "000000000000";
      when "000000000101101" => color_data <= "000000000000";
      when "000000000101110" => color_data <= "000000000000";
      when "000000000101111" => color_data <= "000000000000";
      when "000000000110000" => color_data <= "000000000000";
      when "000000000110001" => color_data <= "000000000000";
      when "000000000110010" => color_data <= "000000000000";
      when "000000000110011" => color_data <= "000000000000";
      when "000000000110100" => color_data <= "000000000000";
      when "000000000110101" => color_data <= "000000000000";
      when "000000000110110" => color_data <= "000000000000";
      when "000000000110111" => color_data <= "000000000000";
      when "000000000111000" => color_data <= "000000000000";
      when "000000000111001" => color_data <= "000000000000";
      when "000000000111010" => color_data <= "000000000000";
      when "000000000111011" => color_data <= "000000000000";
      when "000000000111100" => color_data <= "000000000000";
      when "000000000111101" => color_data <= "000000000000";
      when "000000000111110" => color_data <= "000000000000";
      when "000000000111111" => color_data <= "000000000000";
      when "000000001000000" => color_data <= "000000000000";
      when "000000001000001" => color_data <= "000000000000";
      when "000000001000010" => color_data <= "000000000000";
      when "000000001000011" => color_data <= "000000000000";
      when "000000001000100" => color_data <= "000000000000";
      when "000000001000101" => color_data <= "000000000000";
      when "000000001000110" => color_data <= "000000000000";
      when "000000001000111" => color_data <= "000000000000";
      when "000000001001000" => color_data <= "000000000000";
      when "000000001001001" => color_data <= "000000000000";
      when "000000001001010" => color_data <= "000000000000";
      when "000000001001011" => color_data <= "000000000000";
      when "000000001001100" => color_data <= "000000000000";
      when "000000001001101" => color_data <= "000000000000";
      when "000000001001110" => color_data <= "000000000000";
      when "000000001001111" => color_data <= "000000000000";
      when "000000001010000" => color_data <= "000000000000";
      when "000000001010001" => color_data <= "000000000000";
      when "000000001010010" => color_data <= "000000000000";
      when "000000001010011" => color_data <= "000000000000";
      when "000000001010100" => color_data <= "000000000000";
      when "000000001010101" => color_data <= "000000000000";
      when "000000001010110" => color_data <= "000000000000";
      when "000000001010111" => color_data <= "000000000000";
      when "000000001011000" => color_data <= "000000000000";
      when "000000001011001" => color_data <= "000000000000";
      when "000000001011010" => color_data <= "000000000000";
      when "000000001011011" => color_data <= "000000000000";
      when "000000001011100" => color_data <= "000000000000";
      when "000000001011101" => color_data <= "000000000000";
      when "000000001011110" => color_data <= "000000000000";
      when "000000001011111" => color_data <= "000000000000";
      when "000000001100000" => color_data <= "000000000000";
      when "000000001100001" => color_data <= "000000000000";
      when "000000001100010" => color_data <= "000000000000";
      when "000000001100011" => color_data <= "000000000000";
      when "000000010000000" => color_data <= "000000000000";
      when "000000010000001" => color_data <= "000000000000";
      when "000000010000010" => color_data <= "000000000000";
      when "000000010000011" => color_data <= "000000000000";
      when "000000010000100" => color_data <= "000000000000";
      when "000000010000101" => color_data <= "000000000000";
      when "000000010000110" => color_data <= "000000000000";
      when "000000010000111" => color_data <= "000000000000";
      when "000000010001000" => color_data <= "000000000000";
      when "000000010001001" => color_data <= "000000000000";
      when "000000010001010" => color_data <= "000000000000";
      when "000000010001011" => color_data <= "000000000000";
      when "000000010001100" => color_data <= "000000000000";
      when "000000010001101" => color_data <= "000000000000";
      when "000000010001110" => color_data <= "000000000000";
      when "000000010001111" => color_data <= "000000000000";
      when "000000010010000" => color_data <= "000000000000";
      when "000000010010001" => color_data <= "000000000000";
      when "000000010010010" => color_data <= "000000000000";
      when "000000010010011" => color_data <= "000000000000";
      when "000000010010100" => color_data <= "000000000000";
      when "000000010010101" => color_data <= "000000000000";
      when "000000010010110" => color_data <= "000000000000";
      when "000000010010111" => color_data <= "000000000000";
      when "000000010011000" => color_data <= "000000000000";
      when "000000010011001" => color_data <= "000000000000";
      when "000000010011010" => color_data <= "000000000000";
      when "000000010011011" => color_data <= "000000000000";
      when "000000010011100" => color_data <= "000000000000";
      when "000000010011101" => color_data <= "000000000000";
      when "000000010011110" => color_data <= "000000000000";
      when "000000010011111" => color_data <= "000000000000";
      when "000000010100000" => color_data <= "000000000000";
      when "000000010100001" => color_data <= "000000000000";
      when "000000010100010" => color_data <= "000000000000";
      when "000000010100011" => color_data <= "000000000000";
      when "000000010100100" => color_data <= "000000000000";
      when "000000010100101" => color_data <= "000000000000";
      when "000000010100110" => color_data <= "000000000000";
      when "000000010100111" => color_data <= "000000000000";
      when "000000010101000" => color_data <= "000000000000";
      when "000000010101001" => color_data <= "000000000000";
      when "000000010101010" => color_data <= "000000000000";
      when "000000010101011" => color_data <= "000000000000";
      when "000000010101100" => color_data <= "000000000000";
      when "000000010101101" => color_data <= "000000000000";
      when "000000010101110" => color_data <= "000000000000";
      when "000000010101111" => color_data <= "000000000000";
      when "000000010110000" => color_data <= "000000000000";
      when "000000010110001" => color_data <= "000000000000";
      when "000000010110010" => color_data <= "000000000000";
      when "000000010110011" => color_data <= "000000000000";
      when "000000010110100" => color_data <= "000000000000";
      when "000000010110101" => color_data <= "000000000000";
      when "000000010110110" => color_data <= "000000000000";
      when "000000010110111" => color_data <= "000000000000";
      when "000000010111000" => color_data <= "000000000000";
      when "000000010111001" => color_data <= "000000000000";
      when "000000010111010" => color_data <= "000000000000";
      when "000000010111011" => color_data <= "000000000000";
      when "000000010111100" => color_data <= "000000000000";
      when "000000010111101" => color_data <= "000000000000";
      when "000000010111110" => color_data <= "000000000000";
      when "000000010111111" => color_data <= "000000000000";
      when "000000011000000" => color_data <= "000000000000";
      when "000000011000001" => color_data <= "000000000000";
      when "000000011000010" => color_data <= "000000000000";
      when "000000011000011" => color_data <= "000000000000";
      when "000000011000100" => color_data <= "000000000000";
      when "000000011000101" => color_data <= "000000000000";
      when "000000011000110" => color_data <= "000000000000";
      when "000000011000111" => color_data <= "000000000000";
      when "000000011001000" => color_data <= "000000000000";
      when "000000011001001" => color_data <= "000000000000";
      when "000000011001010" => color_data <= "000000000000";
      when "000000011001011" => color_data <= "000000000000";
      when "000000011001100" => color_data <= "000000000000";
      when "000000011001101" => color_data <= "000000000000";
      when "000000011001110" => color_data <= "000000000000";
      when "000000011001111" => color_data <= "000000000000";
      when "000000011010000" => color_data <= "000000000000";
      when "000000011010001" => color_data <= "000000000000";
      when "000000011010010" => color_data <= "000000000000";
      when "000000011010011" => color_data <= "000000000000";
      when "000000011010100" => color_data <= "000000000000";
      when "000000011010101" => color_data <= "000000000000";
      when "000000011010110" => color_data <= "000000000000";
      when "000000011010111" => color_data <= "000000000000";
      when "000000011011000" => color_data <= "000000000000";
      when "000000011011001" => color_data <= "000000000000";
      when "000000011011010" => color_data <= "000000000000";
      when "000000011011011" => color_data <= "000000000000";
      when "000000011011100" => color_data <= "000000000000";
      when "000000011011101" => color_data <= "000000000000";
      when "000000011011110" => color_data <= "000000000000";
      when "000000011011111" => color_data <= "000000000000";
      when "000000011100000" => color_data <= "000000000000";
      when "000000011100001" => color_data <= "000000000000";
      when "000000011100010" => color_data <= "000000000000";
      when "000000011100011" => color_data <= "000000000000";
      when "000000100000000" => color_data <= "000000000000";
      when "000000100000001" => color_data <= "000000000000";
      when "000000100000010" => color_data <= "000000000000";
      when "000000100000011" => color_data <= "000000000000";
      when "000000100000100" => color_data <= "000000000000";
      when "000000100000101" => color_data <= "000000000000";
      when "000000100000110" => color_data <= "000000000000";
      when "000000100000111" => color_data <= "000000000000";
      when "000000100001000" => color_data <= "000000000000";
      when "000000100001001" => color_data <= "000000000000";
      when "000000100001010" => color_data <= "000000000000";
      when "000000100001011" => color_data <= "000000000000";
      when "000000100001100" => color_data <= "000000000000";
      when "000000100001101" => color_data <= "000000000000";
      when "000000100001110" => color_data <= "000000000000";
      when "000000100001111" => color_data <= "000000000000";
      when "000000100010000" => color_data <= "000000000000";
      when "000000100010001" => color_data <= "000000000000";
      when "000000100010010" => color_data <= "000000000000";
      when "000000100010011" => color_data <= "000000000000";
      when "000000100010100" => color_data <= "000000000000";
      when "000000100010101" => color_data <= "000000000000";
      when "000000100010110" => color_data <= "000000000000";
      when "000000100010111" => color_data <= "000000000000";
      when "000000100011000" => color_data <= "000000000000";
      when "000000100011001" => color_data <= "000000000000";
      when "000000100011010" => color_data <= "000000000000";
      when "000000100011011" => color_data <= "000000000000";
      when "000000100011100" => color_data <= "000000000000";
      when "000000100011101" => color_data <= "000000000000";
      when "000000100011110" => color_data <= "000000000000";
      when "000000100011111" => color_data <= "000000000000";
      when "000000100100000" => color_data <= "000000000000";
      when "000000100100001" => color_data <= "000000000000";
      when "000000100100010" => color_data <= "000000000000";
      when "000000100100011" => color_data <= "000000000000";
      when "000000100100100" => color_data <= "000000000000";
      when "000000100100101" => color_data <= "000000000000";
      when "000000100100110" => color_data <= "000000000000";
      when "000000100100111" => color_data <= "000000000000";
      when "000000100101000" => color_data <= "000000000000";
      when "000000100101001" => color_data <= "000000000000";
      when "000000100101010" => color_data <= "000000000000";
      when "000000100101011" => color_data <= "000000000000";
      when "000000100101100" => color_data <= "000000000000";
      when "000000100101101" => color_data <= "000000000000";
      when "000000100101110" => color_data <= "000000000000";
      when "000000100101111" => color_data <= "000000000000";
      when "000000100110000" => color_data <= "000000000000";
      when "000000100110001" => color_data <= "000000000000";
      when "000000100110010" => color_data <= "000000000000";
      when "000000100110011" => color_data <= "000000000000";
      when "000000100110100" => color_data <= "000000000000";
      when "000000100110101" => color_data <= "000000000000";
      when "000000100110110" => color_data <= "000000000000";
      when "000000100110111" => color_data <= "000000000000";
      when "000000100111000" => color_data <= "000000000000";
      when "000000100111001" => color_data <= "000000000000";
      when "000000100111010" => color_data <= "000000000000";
      when "000000100111011" => color_data <= "000000000000";
      when "000000100111100" => color_data <= "000000000000";
      when "000000100111101" => color_data <= "000000000000";
      when "000000100111110" => color_data <= "000000000000";
      when "000000100111111" => color_data <= "000000000000";
      when "000000101000000" => color_data <= "000000000000";
      when "000000101000001" => color_data <= "000000000000";
      when "000000101000010" => color_data <= "000000000000";
      when "000000101000011" => color_data <= "000000000000";
      when "000000101000100" => color_data <= "000000000000";
      when "000000101000101" => color_data <= "000000000000";
      when "000000101000110" => color_data <= "000000000000";
      when "000000101000111" => color_data <= "000000000000";
      when "000000101001000" => color_data <= "000000000000";
      when "000000101001001" => color_data <= "000000000000";
      when "000000101001010" => color_data <= "000000000000";
      when "000000101001011" => color_data <= "000000000000";
      when "000000101001100" => color_data <= "000000000000";
      when "000000101001101" => color_data <= "000000000000";
      when "000000101001110" => color_data <= "000000000000";
      when "000000101001111" => color_data <= "000000000000";
      when "000000101010000" => color_data <= "000000000000";
      when "000000101010001" => color_data <= "000000000000";
      when "000000101010010" => color_data <= "000000000000";
      when "000000101010011" => color_data <= "000000000000";
      when "000000101010100" => color_data <= "000000000000";
      when "000000101010101" => color_data <= "000000000000";
      when "000000101010110" => color_data <= "000000000000";
      when "000000101010111" => color_data <= "000000000000";
      when "000000101011000" => color_data <= "000000000000";
      when "000000101011001" => color_data <= "000000000000";
      when "000000101011010" => color_data <= "000000000000";
      when "000000101011011" => color_data <= "000000000000";
      when "000000101011100" => color_data <= "000000000000";
      when "000000101011101" => color_data <= "000000000000";
      when "000000101011110" => color_data <= "000000000000";
      when "000000101011111" => color_data <= "000000000000";
      when "000000101100000" => color_data <= "000000000000";
      when "000000101100001" => color_data <= "000000000000";
      when "000000101100010" => color_data <= "000000000000";
      when "000000101100011" => color_data <= "000000000000";
      when "000000110000000" => color_data <= "000000000000";
      when "000000110000001" => color_data <= "000000000000";
      when "000000110000010" => color_data <= "000000000000";
      when "000000110000011" => color_data <= "000000000000";
      when "000000110000100" => color_data <= "000000000000";
      when "000000110000101" => color_data <= "000000000000";
      when "000000110000110" => color_data <= "000000000000";
      when "000000110000111" => color_data <= "000000000000";
      when "000000110001000" => color_data <= "000000000000";
      when "000000110001001" => color_data <= "000000000000";
      when "000000110001010" => color_data <= "000000000000";
      when "000000110001011" => color_data <= "000000000000";
      when "000000110001100" => color_data <= "000000000000";
      when "000000110001101" => color_data <= "000000000000";
      when "000000110001110" => color_data <= "000000000000";
      when "000000110001111" => color_data <= "000000000000";
      when "000000110010000" => color_data <= "000000000000";
      when "000000110010001" => color_data <= "000000000000";
      when "000000110010010" => color_data <= "000000000000";
      when "000000110010011" => color_data <= "000000000000";
      when "000000110010100" => color_data <= "000000000000";
      when "000000110010101" => color_data <= "000000000000";
      when "000000110010110" => color_data <= "000000000000";
      when "000000110010111" => color_data <= "000000000000";
      when "000000110011000" => color_data <= "000000000000";
      when "000000110011001" => color_data <= "000000000000";
      when "000000110011010" => color_data <= "000000000000";
      when "000000110011011" => color_data <= "000000000000";
      when "000000110011100" => color_data <= "000000000000";
      when "000000110011101" => color_data <= "000000000000";
      when "000000110011110" => color_data <= "000000000000";
      when "000000110011111" => color_data <= "000000000000";
      when "000000110100000" => color_data <= "000000000000";
      when "000000110100001" => color_data <= "000000000000";
      when "000000110100010" => color_data <= "000000000000";
      when "000000110100011" => color_data <= "000000000000";
      when "000000110100100" => color_data <= "000000000000";
      when "000000110100101" => color_data <= "000000000000";
      when "000000110100110" => color_data <= "000000000000";
      when "000000110100111" => color_data <= "000000000000";
      when "000000110101000" => color_data <= "000000000000";
      when "000000110101001" => color_data <= "000000000000";
      when "000000110101010" => color_data <= "000000000000";
      when "000000110101011" => color_data <= "000000000000";
      when "000000110101100" => color_data <= "000000000000";
      when "000000110101101" => color_data <= "000000000000";
      when "000000110101110" => color_data <= "000000000000";
      when "000000110101111" => color_data <= "000000000000";
      when "000000110110000" => color_data <= "000000000000";
      when "000000110110001" => color_data <= "000000000000";
      when "000000110110010" => color_data <= "000000000000";
      when "000000110110011" => color_data <= "000000000000";
      when "000000110110100" => color_data <= "000000000000";
      when "000000110110101" => color_data <= "000000000000";
      when "000000110110110" => color_data <= "000000000000";
      when "000000110110111" => color_data <= "000000000000";
      when "000000110111000" => color_data <= "000000000000";
      when "000000110111001" => color_data <= "000000000000";
      when "000000110111010" => color_data <= "000000000000";
      when "000000110111011" => color_data <= "000000000000";
      when "000000110111100" => color_data <= "000000000000";
      when "000000110111101" => color_data <= "000000000000";
      when "000000110111110" => color_data <= "000000000000";
      when "000000110111111" => color_data <= "000000000000";
      when "000000111000000" => color_data <= "000000000000";
      when "000000111000001" => color_data <= "000000000000";
      when "000000111000010" => color_data <= "000000000000";
      when "000000111000011" => color_data <= "000000000000";
      when "000000111000100" => color_data <= "000000000000";
      when "000000111000101" => color_data <= "000000000000";
      when "000000111000110" => color_data <= "000000000000";
      when "000000111000111" => color_data <= "000000000000";
      when "000000111001000" => color_data <= "000000000000";
      when "000000111001001" => color_data <= "000000000000";
      when "000000111001010" => color_data <= "000000000000";
      when "000000111001011" => color_data <= "000000000000";
      when "000000111001100" => color_data <= "000000000000";
      when "000000111001101" => color_data <= "000000000000";
      when "000000111001110" => color_data <= "000000000000";
      when "000000111001111" => color_data <= "000000000000";
      when "000000111010000" => color_data <= "000000000000";
      when "000000111010001" => color_data <= "000000000000";
      when "000000111010010" => color_data <= "000000000000";
      when "000000111010011" => color_data <= "000000000000";
      when "000000111010100" => color_data <= "000000000000";
      when "000000111010101" => color_data <= "000000000000";
      when "000000111010110" => color_data <= "000000000000";
      when "000000111010111" => color_data <= "000000000000";
      when "000000111011000" => color_data <= "000000000000";
      when "000000111011001" => color_data <= "000000000000";
      when "000000111011010" => color_data <= "000000000000";
      when "000000111011011" => color_data <= "000000000000";
      when "000000111011100" => color_data <= "000000000000";
      when "000000111011101" => color_data <= "000000000000";
      when "000000111011110" => color_data <= "000000000000";
      when "000000111011111" => color_data <= "000000000000";
      when "000000111100000" => color_data <= "000000000000";
      when "000000111100001" => color_data <= "000000000000";
      when "000000111100010" => color_data <= "000000000000";
      when "000000111100011" => color_data <= "000000000000";
      when "000001000000000" => color_data <= "000000000000";
      when "000001000000001" => color_data <= "000000000000";
      when "000001000000010" => color_data <= "000000000000";
      when "000001000000011" => color_data <= "000000000000";
      when "000001000000100" => color_data <= "000000000000";
      when "000001000000101" => color_data <= "000000000000";
      when "000001000000110" => color_data <= "000000000000";
      when "000001000000111" => color_data <= "000000000000";
      when "000001000001000" => color_data <= "000000000000";
      when "000001000001001" => color_data <= "000000000000";
      when "000001000001010" => color_data <= "000000000000";
      when "000001000001011" => color_data <= "000000000000";
      when "000001000001100" => color_data <= "000000000000";
      when "000001000001101" => color_data <= "000000000000";
      when "000001000001110" => color_data <= "000000000000";
      when "000001000001111" => color_data <= "000000000000";
      when "000001000010000" => color_data <= "000000000000";
      when "000001000010001" => color_data <= "000000000000";
      when "000001000010010" => color_data <= "000000000000";
      when "000001000010011" => color_data <= "000000000000";
      when "000001000010100" => color_data <= "000000000000";
      when "000001000010101" => color_data <= "000000000000";
      when "000001000010110" => color_data <= "000000000000";
      when "000001000010111" => color_data <= "000000000000";
      when "000001000011000" => color_data <= "000000000000";
      when "000001000011001" => color_data <= "000000000000";
      when "000001000011010" => color_data <= "000000000000";
      when "000001000011011" => color_data <= "000000000000";
      when "000001000011100" => color_data <= "000000000000";
      when "000001000011101" => color_data <= "000000000000";
      when "000001000011110" => color_data <= "000000000000";
      when "000001000011111" => color_data <= "000000000000";
      when "000001000100000" => color_data <= "000000000000";
      when "000001000100001" => color_data <= "000000000000";
      when "000001000100010" => color_data <= "000000000000";
      when "000001000100011" => color_data <= "000000000000";
      when "000001000100100" => color_data <= "000000000000";
      when "000001000100101" => color_data <= "000000000000";
      when "000001000100110" => color_data <= "000000000000";
      when "000001000100111" => color_data <= "000000000000";
      when "000001000101000" => color_data <= "000000000000";
      when "000001000101001" => color_data <= "000000000000";
      when "000001000101010" => color_data <= "000000000000";
      when "000001000101011" => color_data <= "000000000000";
      when "000001000101100" => color_data <= "000000000000";
      when "000001000101101" => color_data <= "000000000000";
      when "000001000101110" => color_data <= "000000000000";
      when "000001000101111" => color_data <= "000000000000";
      when "000001000110000" => color_data <= "000000000000";
      when "000001000110001" => color_data <= "000000000000";
      when "000001000110010" => color_data <= "000000000000";
      when "000001000110011" => color_data <= "000000000000";
      when "000001000110100" => color_data <= "000000000000";
      when "000001000110101" => color_data <= "000000000000";
      when "000001000110110" => color_data <= "000000000000";
      when "000001000110111" => color_data <= "000000000000";
      when "000001000111000" => color_data <= "000000000000";
      when "000001000111001" => color_data <= "000000000000";
      when "000001000111010" => color_data <= "000000000000";
      when "000001000111011" => color_data <= "000000000000";
      when "000001000111100" => color_data <= "000000000000";
      when "000001000111101" => color_data <= "000000000000";
      when "000001000111110" => color_data <= "000000000000";
      when "000001000111111" => color_data <= "000000000000";
      when "000001001000000" => color_data <= "000000000000";
      when "000001001000001" => color_data <= "000000000000";
      when "000001001000010" => color_data <= "000000000000";
      when "000001001000011" => color_data <= "000000000000";
      when "000001001000100" => color_data <= "000000000000";
      when "000001001000101" => color_data <= "000000000000";
      when "000001001000110" => color_data <= "000000000000";
      when "000001001000111" => color_data <= "000000000000";
      when "000001001001000" => color_data <= "000000000000";
      when "000001001001001" => color_data <= "000000000000";
      when "000001001001010" => color_data <= "000000000000";
      when "000001001001011" => color_data <= "000000000000";
      when "000001001001100" => color_data <= "000000000000";
      when "000001001001101" => color_data <= "000000000000";
      when "000001001001110" => color_data <= "000000000000";
      when "000001001001111" => color_data <= "000000000000";
      when "000001001010000" => color_data <= "000000000000";
      when "000001001010001" => color_data <= "000000000000";
      when "000001001010010" => color_data <= "000000000000";
      when "000001001010011" => color_data <= "000000000000";
      when "000001001010100" => color_data <= "000000000000";
      when "000001001010101" => color_data <= "000000000000";
      when "000001001010110" => color_data <= "000000000000";
      when "000001001010111" => color_data <= "000000000000";
      when "000001001011000" => color_data <= "000000000000";
      when "000001001011001" => color_data <= "000000000000";
      when "000001001011010" => color_data <= "000000000000";
      when "000001001011011" => color_data <= "000000000000";
      when "000001001011100" => color_data <= "000000000000";
      when "000001001011101" => color_data <= "000000000000";
      when "000001001011110" => color_data <= "000000000000";
      when "000001001011111" => color_data <= "000000000000";
      when "000001001100000" => color_data <= "000000000000";
      when "000001001100001" => color_data <= "000000000000";
      when "000001001100010" => color_data <= "000000000000";
      when "000001001100011" => color_data <= "000000000000";
      when "000001010000000" => color_data <= "000000000000";
      when "000001010000001" => color_data <= "000000000000";
      when "000001010000010" => color_data <= "000000000000";
      when "000001010000011" => color_data <= "000000000000";
      when "000001010000100" => color_data <= "000000000000";
      when "000001010000101" => color_data <= "000000000000";
      when "000001010000110" => color_data <= "000000000000";
      when "000001010000111" => color_data <= "000000000000";
      when "000001010001000" => color_data <= "000000000000";
      when "000001010001001" => color_data <= "000000000000";
      when "000001010001010" => color_data <= "000000000000";
      when "000001010001011" => color_data <= "000000000000";
      when "000001010001100" => color_data <= "000000000000";
      when "000001010001101" => color_data <= "000000000000";
      when "000001010001110" => color_data <= "000000000000";
      when "000001010001111" => color_data <= "000000000000";
      when "000001010010000" => color_data <= "000000000000";
      when "000001010010001" => color_data <= "000000000000";
      when "000001010010010" => color_data <= "000000000000";
      when "000001010010011" => color_data <= "000000000000";
      when "000001010010100" => color_data <= "000000000000";
      when "000001010010101" => color_data <= "000000000000";
      when "000001010010110" => color_data <= "000000000000";
      when "000001010010111" => color_data <= "000000000000";
      when "000001010011000" => color_data <= "000000000000";
      when "000001010011001" => color_data <= "000000000000";
      when "000001010011010" => color_data <= "000000000000";
      when "000001010011011" => color_data <= "000000000000";
      when "000001010011100" => color_data <= "000000000000";
      when "000001010011101" => color_data <= "000000000000";
      when "000001010011110" => color_data <= "000000000000";
      when "000001010011111" => color_data <= "000000000000";
      when "000001010100000" => color_data <= "000000000000";
      when "000001010100001" => color_data <= "000000000000";
      when "000001010100010" => color_data <= "000000000000";
      when "000001010100011" => color_data <= "000000000000";
      when "000001010100100" => color_data <= "000000000000";
      when "000001010100101" => color_data <= "000000000000";
      when "000001010100110" => color_data <= "000000000000";
      when "000001010100111" => color_data <= "000000000000";
      when "000001010101000" => color_data <= "000000000000";
      when "000001010101001" => color_data <= "000000000000";
      when "000001010101010" => color_data <= "000000000000";
      when "000001010101011" => color_data <= "000000000000";
      when "000001010101100" => color_data <= "000000000000";
      when "000001010101101" => color_data <= "000000000000";
      when "000001010101110" => color_data <= "000000000000";
      when "000001010101111" => color_data <= "000000000000";
      when "000001010110000" => color_data <= "000000000000";
      when "000001010110001" => color_data <= "000000000000";
      when "000001010110010" => color_data <= "000000000000";
      when "000001010110011" => color_data <= "000000000000";
      when "000001010110100" => color_data <= "000000000000";
      when "000001010110101" => color_data <= "000000000000";
      when "000001010110110" => color_data <= "000000000000";
      when "000001010110111" => color_data <= "000000000000";
      when "000001010111000" => color_data <= "000000000000";
      when "000001010111001" => color_data <= "000000000000";
      when "000001010111010" => color_data <= "000000000000";
      when "000001010111011" => color_data <= "000000000000";
      when "000001010111100" => color_data <= "000000000000";
      when "000001010111101" => color_data <= "000000000000";
      when "000001010111110" => color_data <= "000000000000";
      when "000001010111111" => color_data <= "000000000000";
      when "000001011000000" => color_data <= "000000000000";
      when "000001011000001" => color_data <= "000000000000";
      when "000001011000010" => color_data <= "000000000000";
      when "000001011000011" => color_data <= "000000000000";
      when "000001011000100" => color_data <= "000000000000";
      when "000001011000101" => color_data <= "000000000000";
      when "000001011000110" => color_data <= "000000000000";
      when "000001011000111" => color_data <= "000000000000";
      when "000001011001000" => color_data <= "000000000000";
      when "000001011001001" => color_data <= "000000000000";
      when "000001011001010" => color_data <= "000000000000";
      when "000001011001011" => color_data <= "000000000000";
      when "000001011001100" => color_data <= "000000000000";
      when "000001011001101" => color_data <= "000000000000";
      when "000001011001110" => color_data <= "000000000000";
      when "000001011001111" => color_data <= "000000000000";
      when "000001011010000" => color_data <= "000000000000";
      when "000001011010001" => color_data <= "000000000000";
      when "000001011010010" => color_data <= "000000000000";
      when "000001011010011" => color_data <= "000000000000";
      when "000001011010100" => color_data <= "000000000000";
      when "000001011010101" => color_data <= "000000000000";
      when "000001011010110" => color_data <= "000000000000";
      when "000001011010111" => color_data <= "000000000000";
      when "000001011011000" => color_data <= "000000000000";
      when "000001011011001" => color_data <= "000000000000";
      when "000001011011010" => color_data <= "000000000000";
      when "000001011011011" => color_data <= "000000000000";
      when "000001011011100" => color_data <= "000000000000";
      when "000001011011101" => color_data <= "000000000000";
      when "000001011011110" => color_data <= "000000000000";
      when "000001011011111" => color_data <= "000000000000";
      when "000001011100000" => color_data <= "000000000000";
      when "000001011100001" => color_data <= "000000000000";
      when "000001011100010" => color_data <= "000000000000";
      when "000001011100011" => color_data <= "000000000000";
      when "000001100000000" => color_data <= "000000000000";
      when "000001100000001" => color_data <= "000000000000";
      when "000001100000010" => color_data <= "000000000000";
      when "000001100000011" => color_data <= "000000000000";
      when "000001100000100" => color_data <= "000000000000";
      when "000001100000101" => color_data <= "000000000000";
      when "000001100000110" => color_data <= "000000000000";
      when "000001100000111" => color_data <= "000000000000";
      when "000001100001000" => color_data <= "000000000000";
      when "000001100001001" => color_data <= "000000000000";
      when "000001100001010" => color_data <= "000000000000";
      when "000001100001011" => color_data <= "000000000000";
      when "000001100001100" => color_data <= "000000000000";
      when "000001100001101" => color_data <= "000000000000";
      when "000001100001110" => color_data <= "000000000000";
      when "000001100001111" => color_data <= "000000000000";
      when "000001100010000" => color_data <= "000000000000";
      when "000001100010001" => color_data <= "000000000000";
      when "000001100010010" => color_data <= "000000000000";
      when "000001100010011" => color_data <= "000000000000";
      when "000001100010100" => color_data <= "000000000000";
      when "000001100010101" => color_data <= "000000000000";
      when "000001100010110" => color_data <= "000000000000";
      when "000001100010111" => color_data <= "000000000000";
      when "000001100011000" => color_data <= "000000000000";
      when "000001100011001" => color_data <= "000000000000";
      when "000001100011010" => color_data <= "000000000000";
      when "000001100011011" => color_data <= "000000000000";
      when "000001100011100" => color_data <= "000000000000";
      when "000001100011101" => color_data <= "000000000000";
      when "000001100011110" => color_data <= "000000000000";
      when "000001100011111" => color_data <= "000000000000";
      when "000001100100000" => color_data <= "000000000000";
      when "000001100100001" => color_data <= "000000000000";
      when "000001100100010" => color_data <= "000000000000";
      when "000001100100011" => color_data <= "000000000000";
      when "000001100100100" => color_data <= "000000000000";
      when "000001100100101" => color_data <= "000000000000";
      when "000001100100110" => color_data <= "000000000000";
      when "000001100100111" => color_data <= "000000000000";
      when "000001100101000" => color_data <= "000000000000";
      when "000001100101001" => color_data <= "000000000000";
      when "000001100101010" => color_data <= "000000000000";
      when "000001100101011" => color_data <= "000000000000";
      when "000001100101100" => color_data <= "000000000000";
      when "000001100101101" => color_data <= "000000000000";
      when "000001100101110" => color_data <= "000000000000";
      when "000001100101111" => color_data <= "000000000000";
      when "000001100110000" => color_data <= "000000000000";
      when "000001100110001" => color_data <= "000000000000";
      when "000001100110010" => color_data <= "000000000000";
      when "000001100110011" => color_data <= "000000000000";
      when "000001100110100" => color_data <= "000000000000";
      when "000001100110101" => color_data <= "000000000000";
      when "000001100110110" => color_data <= "000000000000";
      when "000001100110111" => color_data <= "000000000000";
      when "000001100111000" => color_data <= "000000000000";
      when "000001100111001" => color_data <= "000000000000";
      when "000001100111010" => color_data <= "000000000000";
      when "000001100111011" => color_data <= "000000000000";
      when "000001100111100" => color_data <= "000000000000";
      when "000001100111101" => color_data <= "000000000000";
      when "000001100111110" => color_data <= "000000000000";
      when "000001100111111" => color_data <= "000000000000";
      when "000001101000000" => color_data <= "000000000000";
      when "000001101000001" => color_data <= "000000000000";
      when "000001101000010" => color_data <= "000000000000";
      when "000001101000011" => color_data <= "000000000000";
      when "000001101000100" => color_data <= "000000000000";
      when "000001101000101" => color_data <= "000000000000";
      when "000001101000110" => color_data <= "000000000000";
      when "000001101000111" => color_data <= "000000000000";
      when "000001101001000" => color_data <= "000000000000";
      when "000001101001001" => color_data <= "000000000000";
      when "000001101001010" => color_data <= "000000000000";
      when "000001101001011" => color_data <= "000000000000";
      when "000001101001100" => color_data <= "000000000000";
      when "000001101001101" => color_data <= "000000000000";
      when "000001101001110" => color_data <= "000000000000";
      when "000001101001111" => color_data <= "000000000000";
      when "000001101010000" => color_data <= "000000000000";
      when "000001101010001" => color_data <= "000000000000";
      when "000001101010010" => color_data <= "000000000000";
      when "000001101010011" => color_data <= "000000000000";
      when "000001101010100" => color_data <= "000000000000";
      when "000001101010101" => color_data <= "000000000000";
      when "000001101010110" => color_data <= "000000000000";
      when "000001101010111" => color_data <= "000000000000";
      when "000001101011000" => color_data <= "000000000000";
      when "000001101011001" => color_data <= "000000000000";
      when "000001101011010" => color_data <= "000000000000";
      when "000001101011011" => color_data <= "000000000000";
      when "000001101011100" => color_data <= "000000000000";
      when "000001101011101" => color_data <= "000000000000";
      when "000001101011110" => color_data <= "000000000000";
      when "000001101011111" => color_data <= "000000000000";
      when "000001101100000" => color_data <= "000000000000";
      when "000001101100001" => color_data <= "000000000000";
      when "000001101100010" => color_data <= "000000000000";
      when "000001101100011" => color_data <= "000000000000";
      when "000001110000000" => color_data <= "000000000000";
      when "000001110000001" => color_data <= "000000000000";
      when "000001110000010" => color_data <= "000000000000";
      when "000001110000011" => color_data <= "000000000000";
      when "000001110000100" => color_data <= "000000000000";
      when "000001110000101" => color_data <= "000000000000";
      when "000001110000110" => color_data <= "000000000000";
      when "000001110000111" => color_data <= "000000000000";
      when "000001110001000" => color_data <= "000000000000";
      when "000001110001001" => color_data <= "000000000000";
      when "000001110001010" => color_data <= "000000000000";
      when "000001110001011" => color_data <= "000000000000";
      when "000001110001100" => color_data <= "000000000000";
      when "000001110001101" => color_data <= "000000000000";
      when "000001110001110" => color_data <= "000000000000";
      when "000001110001111" => color_data <= "000000000000";
      when "000001110010000" => color_data <= "000000000000";
      when "000001110010001" => color_data <= "000000000000";
      when "000001110010010" => color_data <= "000000000000";
      when "000001110010011" => color_data <= "000000000000";
      when "000001110010100" => color_data <= "000000000000";
      when "000001110010101" => color_data <= "000000000000";
      when "000001110010110" => color_data <= "000000000000";
      when "000001110010111" => color_data <= "000000000000";
      when "000001110011000" => color_data <= "000000000000";
      when "000001110011001" => color_data <= "000000000000";
      when "000001110011010" => color_data <= "000000000000";
      when "000001110011011" => color_data <= "000000000000";
      when "000001110011100" => color_data <= "000000000000";
      when "000001110011101" => color_data <= "000000000000";
      when "000001110011110" => color_data <= "000000000000";
      when "000001110011111" => color_data <= "000000000000";
      when "000001110100000" => color_data <= "000000000000";
      when "000001110100001" => color_data <= "000000000000";
      when "000001110100010" => color_data <= "000000000000";
      when "000001110100011" => color_data <= "000000000000";
      when "000001110100100" => color_data <= "000000000000";
      when "000001110100101" => color_data <= "000000000000";
      when "000001110100110" => color_data <= "000000000000";
      when "000001110100111" => color_data <= "000000000000";
      when "000001110101000" => color_data <= "000000000000";
      when "000001110101001" => color_data <= "000000000000";
      when "000001110101010" => color_data <= "000000000000";
      when "000001110101011" => color_data <= "000000000000";
      when "000001110101100" => color_data <= "000000000000";
      when "000001110101101" => color_data <= "000000000000";
      when "000001110101110" => color_data <= "000000000000";
      when "000001110101111" => color_data <= "000000000000";
      when "000001110110000" => color_data <= "000000000000";
      when "000001110110001" => color_data <= "000000000000";
      when "000001110110010" => color_data <= "000000000000";
      when "000001110110011" => color_data <= "000000000000";
      when "000001110110100" => color_data <= "000000000000";
      when "000001110110101" => color_data <= "000000000000";
      when "000001110110110" => color_data <= "000000000000";
      when "000001110110111" => color_data <= "000000000000";
      when "000001110111000" => color_data <= "000000000000";
      when "000001110111001" => color_data <= "000000000000";
      when "000001110111010" => color_data <= "000000000000";
      when "000001110111011" => color_data <= "000000000000";
      when "000001110111100" => color_data <= "000000000000";
      when "000001110111101" => color_data <= "000000000000";
      when "000001110111110" => color_data <= "000000000000";
      when "000001110111111" => color_data <= "000000000000";
      when "000001111000000" => color_data <= "000000000000";
      when "000001111000001" => color_data <= "000000000000";
      when "000001111000010" => color_data <= "000000000000";
      when "000001111000011" => color_data <= "000000000000";
      when "000001111000100" => color_data <= "000000000000";
      when "000001111000101" => color_data <= "000000000000";
      when "000001111000110" => color_data <= "000000000000";
      when "000001111000111" => color_data <= "000000000000";
      when "000001111001000" => color_data <= "000000000000";
      when "000001111001001" => color_data <= "000000000000";
      when "000001111001010" => color_data <= "000000000000";
      when "000001111001011" => color_data <= "000000000000";
      when "000001111001100" => color_data <= "000000000000";
      when "000001111001101" => color_data <= "000000000000";
      when "000001111001110" => color_data <= "000000000000";
      when "000001111001111" => color_data <= "000000000000";
      when "000001111010000" => color_data <= "000000000000";
      when "000001111010001" => color_data <= "000000000000";
      when "000001111010010" => color_data <= "000000000000";
      when "000001111010011" => color_data <= "000000000000";
      when "000001111010100" => color_data <= "000000000000";
      when "000001111010101" => color_data <= "000000000000";
      when "000001111010110" => color_data <= "000000000000";
      when "000001111010111" => color_data <= "000000000000";
      when "000001111011000" => color_data <= "000000000000";
      when "000001111011001" => color_data <= "000000000000";
      when "000001111011010" => color_data <= "000000000000";
      when "000001111011011" => color_data <= "000000000000";
      when "000001111011100" => color_data <= "000000000000";
      when "000001111011101" => color_data <= "000000000000";
      when "000001111011110" => color_data <= "000000000000";
      when "000001111011111" => color_data <= "000000000000";
      when "000001111100000" => color_data <= "000000000000";
      when "000001111100001" => color_data <= "000000000000";
      when "000001111100010" => color_data <= "000000000000";
      when "000001111100011" => color_data <= "000000000000";
      when "000010000000000" => color_data <= "000000000000";
      when "000010000000001" => color_data <= "000000000000";
      when "000010000000010" => color_data <= "000000000000";
      when "000010000000011" => color_data <= "000000000000";
      when "000010000000100" => color_data <= "000000000000";
      when "000010000000101" => color_data <= "000000000000";
      when "000010000000110" => color_data <= "000000000000";
      when "000010000000111" => color_data <= "000000000000";
      when "000010000001000" => color_data <= "000000000000";
      when "000010000001001" => color_data <= "000000000000";
      when "000010000001010" => color_data <= "000000000000";
      when "000010000001011" => color_data <= "000000000000";
      when "000010000001100" => color_data <= "000000000000";
      when "000010000001101" => color_data <= "000000000000";
      when "000010000001110" => color_data <= "000000000000";
      when "000010000001111" => color_data <= "000000000000";
      when "000010000010000" => color_data <= "000000000000";
      when "000010000010001" => color_data <= "000000000000";
      when "000010000010010" => color_data <= "000000000000";
      when "000010000010011" => color_data <= "000000000000";
      when "000010000010100" => color_data <= "000000000000";
      when "000010000010101" => color_data <= "000000000000";
      when "000010000010110" => color_data <= "000000000000";
      when "000010000010111" => color_data <= "000000000000";
      when "000010000011000" => color_data <= "000000000000";
      when "000010000011001" => color_data <= "000000000000";
      when "000010000011010" => color_data <= "000000000000";
      when "000010000011011" => color_data <= "000000000000";
      when "000010000011100" => color_data <= "000000000000";
      when "000010000011101" => color_data <= "000000000000";
      when "000010000011110" => color_data <= "000000000000";
      when "000010000011111" => color_data <= "000000000000";
      when "000010000100000" => color_data <= "000000000000";
      when "000010000100001" => color_data <= "000000000000";
      when "000010000100010" => color_data <= "000000000000";
      when "000010000100011" => color_data <= "000000000000";
      when "000010000100100" => color_data <= "000000000000";
      when "000010000100101" => color_data <= "000000000000";
      when "000010000100110" => color_data <= "000000000000";
      when "000010000100111" => color_data <= "000000000000";
      when "000010000101000" => color_data <= "000000000000";
      when "000010000101001" => color_data <= "000000000000";
      when "000010000101010" => color_data <= "000000000000";
      when "000010000101011" => color_data <= "000000000000";
      when "000010000101100" => color_data <= "000000000000";
      when "000010000101101" => color_data <= "000000000000";
      when "000010000101110" => color_data <= "000100010001";
      when "000010000101111" => color_data <= "001000100001";
      when "000010000110000" => color_data <= "001100110010";
      when "000010000110001" => color_data <= "001100110010";
      when "000010000110010" => color_data <= "010001000010";
      when "000010000110011" => color_data <= "010101000010";
      when "000010000110100" => color_data <= "001100110010";
      when "000010000110101" => color_data <= "001000100001";
      when "000010000110110" => color_data <= "000100010000";
      when "000010000110111" => color_data <= "000000000000";
      when "000010000111000" => color_data <= "000000000000";
      when "000010000111001" => color_data <= "000000000000";
      when "000010000111010" => color_data <= "000000000000";
      when "000010000111011" => color_data <= "000000000000";
      when "000010000111100" => color_data <= "000000000000";
      when "000010000111101" => color_data <= "000000000000";
      when "000010000111110" => color_data <= "000000000000";
      when "000010000111111" => color_data <= "000000000000";
      when "000010001000000" => color_data <= "000000000000";
      when "000010001000001" => color_data <= "000000000000";
      when "000010001000010" => color_data <= "000000000000";
      when "000010001000011" => color_data <= "000000000000";
      when "000010001000100" => color_data <= "000000000000";
      when "000010001000101" => color_data <= "000000000000";
      when "000010001000110" => color_data <= "000000000000";
      when "000010001000111" => color_data <= "000000000000";
      when "000010001001000" => color_data <= "000000000000";
      when "000010001001001" => color_data <= "000000000000";
      when "000010001001010" => color_data <= "000000000000";
      when "000010001001011" => color_data <= "000000000000";
      when "000010001001100" => color_data <= "000000000000";
      when "000010001001101" => color_data <= "000000000000";
      when "000010001001110" => color_data <= "000000000000";
      when "000010001001111" => color_data <= "000000000000";
      when "000010001010000" => color_data <= "000000000000";
      when "000010001010001" => color_data <= "000000000000";
      when "000010001010010" => color_data <= "000000000000";
      when "000010001010011" => color_data <= "000000000000";
      when "000010001010100" => color_data <= "000000000000";
      when "000010001010101" => color_data <= "000000000000";
      when "000010001010110" => color_data <= "000000000000";
      when "000010001010111" => color_data <= "000000000000";
      when "000010001011000" => color_data <= "000000000000";
      when "000010001011001" => color_data <= "000000000000";
      when "000010001011010" => color_data <= "000000000000";
      when "000010001011011" => color_data <= "000000000000";
      when "000010001011100" => color_data <= "000000000000";
      when "000010001011101" => color_data <= "000000000000";
      when "000010001011110" => color_data <= "000000000000";
      when "000010001011111" => color_data <= "000000000000";
      when "000010001100000" => color_data <= "000000000000";
      when "000010001100001" => color_data <= "000000000000";
      when "000010001100010" => color_data <= "000000000000";
      when "000010001100011" => color_data <= "000000000000";
      when "000010010000000" => color_data <= "000000000000";
      when "000010010000001" => color_data <= "000000000000";
      when "000010010000010" => color_data <= "000000000000";
      when "000010010000011" => color_data <= "000000000000";
      when "000010010000100" => color_data <= "000000000000";
      when "000010010000101" => color_data <= "000000000000";
      when "000010010000110" => color_data <= "000000000000";
      when "000010010000111" => color_data <= "000000000000";
      when "000010010001000" => color_data <= "000000000000";
      when "000010010001001" => color_data <= "000000000000";
      when "000010010001010" => color_data <= "000000000000";
      when "000010010001011" => color_data <= "000000000000";
      when "000010010001100" => color_data <= "000000000000";
      when "000010010001101" => color_data <= "000000000000";
      when "000010010001110" => color_data <= "000000000000";
      when "000010010001111" => color_data <= "000000000000";
      when "000010010010000" => color_data <= "000000000000";
      when "000010010010001" => color_data <= "000000000000";
      when "000010010010010" => color_data <= "000000000000";
      when "000010010010011" => color_data <= "000000000000";
      when "000010010010100" => color_data <= "000000000000";
      when "000010010010101" => color_data <= "000000000000";
      when "000010010010110" => color_data <= "000000000000";
      when "000010010010111" => color_data <= "000000000000";
      when "000010010011000" => color_data <= "000000000000";
      when "000010010011001" => color_data <= "000000000000";
      when "000010010011010" => color_data <= "000000000000";
      when "000010010011011" => color_data <= "000000000000";
      when "000010010011100" => color_data <= "000000000000";
      when "000010010011101" => color_data <= "000000000000";
      when "000010010011110" => color_data <= "000000000000";
      when "000010010011111" => color_data <= "000000000000";
      when "000010010100000" => color_data <= "000000000000";
      when "000010010100001" => color_data <= "000000000000";
      when "000010010100010" => color_data <= "000000000000";
      when "000010010100011" => color_data <= "000000000000";
      when "000010010100100" => color_data <= "000000000000";
      when "000010010100101" => color_data <= "000000000000";
      when "000010010100110" => color_data <= "000000000000";
      when "000010010100111" => color_data <= "000000000000";
      when "000010010101000" => color_data <= "000000000000";
      when "000010010101001" => color_data <= "000000000000";
      when "000010010101010" => color_data <= "001100110010";
      when "000010010101011" => color_data <= "011101100011";
      when "000010010101100" => color_data <= "100110000010";
      when "000010010101101" => color_data <= "101110100001";
      when "000010010101110" => color_data <= "110110110000";
      when "000010010101111" => color_data <= "111111010000";
      when "000010010110000" => color_data <= "111111000000";
      when "000010010110001" => color_data <= "111111000000";
      when "000010010110010" => color_data <= "111111010000";
      when "000010010110011" => color_data <= "111111010010";
      when "000010010110100" => color_data <= "111111010000";
      when "000010010110101" => color_data <= "111111000000";
      when "000010010110110" => color_data <= "110110110000";
      when "000010010110111" => color_data <= "101110010001";
      when "000010010111000" => color_data <= "100001110010";
      when "000010010111001" => color_data <= "011001010011";
      when "000010010111010" => color_data <= "001000100001";
      when "000010010111011" => color_data <= "000000000000";
      when "000010010111100" => color_data <= "000000000000";
      when "000010010111101" => color_data <= "000000000000";
      when "000010010111110" => color_data <= "000000000000";
      when "000010010111111" => color_data <= "000000000000";
      when "000010011000000" => color_data <= "000000000000";
      when "000010011000001" => color_data <= "000000000000";
      when "000010011000010" => color_data <= "000000000000";
      when "000010011000011" => color_data <= "000000000000";
      when "000010011000100" => color_data <= "000000000000";
      when "000010011000101" => color_data <= "000000000000";
      when "000010011000110" => color_data <= "000000000000";
      when "000010011000111" => color_data <= "000000000000";
      when "000010011001000" => color_data <= "000000000000";
      when "000010011001001" => color_data <= "000000000000";
      when "000010011001010" => color_data <= "000000000000";
      when "000010011001011" => color_data <= "000000000000";
      when "000010011001100" => color_data <= "000000000000";
      when "000010011001101" => color_data <= "000000000000";
      when "000010011001110" => color_data <= "000000000000";
      when "000010011001111" => color_data <= "000000000000";
      when "000010011010000" => color_data <= "000000000000";
      when "000010011010001" => color_data <= "000000000000";
      when "000010011010010" => color_data <= "000000000000";
      when "000010011010011" => color_data <= "000000000000";
      when "000010011010100" => color_data <= "000000000000";
      when "000010011010101" => color_data <= "000000000000";
      when "000010011010110" => color_data <= "000000000000";
      when "000010011010111" => color_data <= "000000000000";
      when "000010011011000" => color_data <= "000000000000";
      when "000010011011001" => color_data <= "000000000000";
      when "000010011011010" => color_data <= "000000000000";
      when "000010011011011" => color_data <= "000000000000";
      when "000010011011100" => color_data <= "000000000000";
      when "000010011011101" => color_data <= "000000000000";
      when "000010011011110" => color_data <= "000000000000";
      when "000010011011111" => color_data <= "000000000000";
      when "000010011100000" => color_data <= "000000000000";
      when "000010011100001" => color_data <= "000000000000";
      when "000010011100010" => color_data <= "000000000000";
      when "000010011100011" => color_data <= "000000000000";
      when "000010100000000" => color_data <= "000000000000";
      when "000010100000001" => color_data <= "000000000000";
      when "000010100000010" => color_data <= "000000000000";
      when "000010100000011" => color_data <= "000000000000";
      when "000010100000100" => color_data <= "000000000000";
      when "000010100000101" => color_data <= "000000000000";
      when "000010100000110" => color_data <= "000000000000";
      when "000010100000111" => color_data <= "000000000000";
      when "000010100001000" => color_data <= "000000000000";
      when "000010100001001" => color_data <= "000000000000";
      when "000010100001010" => color_data <= "000000000000";
      when "000010100001011" => color_data <= "000000000000";
      when "000010100001100" => color_data <= "000000000000";
      when "000010100001101" => color_data <= "000000000000";
      when "000010100001110" => color_data <= "000000000000";
      when "000010100001111" => color_data <= "000000000000";
      when "000010100010000" => color_data <= "000000000000";
      when "000010100010001" => color_data <= "000000000000";
      when "000010100010010" => color_data <= "000000000000";
      when "000010100010011" => color_data <= "000000000000";
      when "000010100010100" => color_data <= "000000000000";
      when "000010100010101" => color_data <= "000000000000";
      when "000010100010110" => color_data <= "000000000000";
      when "000010100010111" => color_data <= "000000000000";
      when "000010100011000" => color_data <= "000000000000";
      when "000010100011001" => color_data <= "000000000000";
      when "000010100011010" => color_data <= "000000000000";
      when "000010100011011" => color_data <= "000000000000";
      when "000010100011100" => color_data <= "000000000000";
      when "000010100011101" => color_data <= "000000000000";
      when "000010100011110" => color_data <= "000000000000";
      when "000010100011111" => color_data <= "000000000000";
      when "000010100100000" => color_data <= "000000000000";
      when "000010100100001" => color_data <= "000000000000";
      when "000010100100010" => color_data <= "000000000000";
      when "000010100100011" => color_data <= "000000000000";
      when "000010100100100" => color_data <= "000000000000";
      when "000010100100101" => color_data <= "000000000000";
      when "000010100100110" => color_data <= "000000000000";
      when "000010100100111" => color_data <= "010000110010";
      when "000010100101000" => color_data <= "010101010010";
      when "000010100101001" => color_data <= "100001110010";
      when "000010100101010" => color_data <= "110110110000";
      when "000010100101011" => color_data <= "111111000000";
      when "000010100101100" => color_data <= "111111000000";
      when "000010100101101" => color_data <= "111111010000";
      when "000010100101110" => color_data <= "111111010000";
      when "000010100101111" => color_data <= "111111010000";
      when "000010100110000" => color_data <= "111111010000";
      when "000010100110001" => color_data <= "111111010000";
      when "000010100110010" => color_data <= "111111010010";
      when "000010100110011" => color_data <= "111111101001";
      when "000010100110100" => color_data <= "111111010011";
      when "000010100110101" => color_data <= "111111010000";
      when "000010100110110" => color_data <= "111111010000";
      when "000010100110111" => color_data <= "111111010000";
      when "000010100111000" => color_data <= "111111000000";
      when "000010100111001" => color_data <= "111111000000";
      when "000010100111010" => color_data <= "110110110000";
      when "000010100111011" => color_data <= "101110100001";
      when "000010100111100" => color_data <= "011001100011";
      when "000010100111101" => color_data <= "001000100001";
      when "000010100111110" => color_data <= "000000000000";
      when "000010100111111" => color_data <= "000000000000";
      when "000010101000000" => color_data <= "000000000000";
      when "000010101000001" => color_data <= "000000000000";
      when "000010101000010" => color_data <= "000000000000";
      when "000010101000011" => color_data <= "000000000000";
      when "000010101000100" => color_data <= "000000000000";
      when "000010101000101" => color_data <= "000000000000";
      when "000010101000110" => color_data <= "000000000000";
      when "000010101000111" => color_data <= "000000000000";
      when "000010101001000" => color_data <= "000000000000";
      when "000010101001001" => color_data <= "000000000000";
      when "000010101001010" => color_data <= "000000000000";
      when "000010101001011" => color_data <= "000000000000";
      when "000010101001100" => color_data <= "000000000000";
      when "000010101001101" => color_data <= "000000000000";
      when "000010101001110" => color_data <= "000000000000";
      when "000010101001111" => color_data <= "000000000000";
      when "000010101010000" => color_data <= "000000000000";
      when "000010101010001" => color_data <= "000000000000";
      when "000010101010010" => color_data <= "000000000000";
      when "000010101010011" => color_data <= "000000000000";
      when "000010101010100" => color_data <= "000000000000";
      when "000010101010101" => color_data <= "000000000000";
      when "000010101010110" => color_data <= "000000000000";
      when "000010101010111" => color_data <= "000000000000";
      when "000010101011000" => color_data <= "000000000000";
      when "000010101011001" => color_data <= "000000000000";
      when "000010101011010" => color_data <= "000000000000";
      when "000010101011011" => color_data <= "000000000000";
      when "000010101011100" => color_data <= "000000000000";
      when "000010101011101" => color_data <= "000000000000";
      when "000010101011110" => color_data <= "000000000000";
      when "000010101011111" => color_data <= "000000000000";
      when "000010101100000" => color_data <= "000000000000";
      when "000010101100001" => color_data <= "000000000000";
      when "000010101100010" => color_data <= "000000000000";
      when "000010101100011" => color_data <= "000000000000";
      when "000010110000000" => color_data <= "000000000000";
      when "000010110000001" => color_data <= "000000000000";
      when "000010110000010" => color_data <= "000000000000";
      when "000010110000011" => color_data <= "000000000000";
      when "000010110000100" => color_data <= "000000000000";
      when "000010110000101" => color_data <= "000000000000";
      when "000010110000110" => color_data <= "000000000000";
      when "000010110000111" => color_data <= "000000000000";
      when "000010110001000" => color_data <= "000000000000";
      when "000010110001001" => color_data <= "000000000000";
      when "000010110001010" => color_data <= "000000000000";
      when "000010110001011" => color_data <= "000000000000";
      when "000010110001100" => color_data <= "000000000000";
      when "000010110001101" => color_data <= "000000000000";
      when "000010110001110" => color_data <= "000000000000";
      when "000010110001111" => color_data <= "000000000000";
      when "000010110010000" => color_data <= "000000000000";
      when "000010110010001" => color_data <= "000000000000";
      when "000010110010010" => color_data <= "000000000000";
      when "000010110010011" => color_data <= "000000000000";
      when "000010110010100" => color_data <= "000000000000";
      when "000010110010101" => color_data <= "000000000000";
      when "000010110010110" => color_data <= "000000000000";
      when "000010110010111" => color_data <= "000000000000";
      when "000010110011000" => color_data <= "000000000000";
      when "000010110011001" => color_data <= "000000000000";
      when "000010110011010" => color_data <= "000000000000";
      when "000010110011011" => color_data <= "000000000000";
      when "000010110011100" => color_data <= "000000000000";
      when "000010110011101" => color_data <= "000000000000";
      when "000010110011110" => color_data <= "000000000000";
      when "000010110011111" => color_data <= "000000000000";
      when "000010110100000" => color_data <= "000000000000";
      when "000010110100001" => color_data <= "000000000000";
      when "000010110100010" => color_data <= "000000000000";
      when "000010110100011" => color_data <= "000000000000";
      when "000010110100100" => color_data <= "000000000000";
      when "000010110100101" => color_data <= "010101000010";
      when "000010110100110" => color_data <= "100001110010";
      when "000010110100111" => color_data <= "100110000010";
      when "000010110101000" => color_data <= "111111100110";
      when "000010110101001" => color_data <= "111111010010";
      when "000010110101010" => color_data <= "111111010000";
      when "000010110101011" => color_data <= "111111010001";
      when "000010110101100" => color_data <= "111111010000";
      when "000010110101101" => color_data <= "111111010000";
      when "000010110101110" => color_data <= "111111010000";
      when "000010110101111" => color_data <= "111111010000";
      when "000010110110000" => color_data <= "111111010000";
      when "000010110110001" => color_data <= "111111010000";
      when "000010110110010" => color_data <= "111111010011";
      when "000010110110011" => color_data <= "111111101010";
      when "000010110110100" => color_data <= "111111010100";
      when "000010110110101" => color_data <= "111111010000";
      when "000010110110110" => color_data <= "111111010001";
      when "000010110110111" => color_data <= "111111010000";
      when "000010110111000" => color_data <= "111111010000";
      when "000010110111001" => color_data <= "111111010001";
      when "000010110111010" => color_data <= "111111010000";
      when "000010110111011" => color_data <= "111111010000";
      when "000010110111100" => color_data <= "111111000000";
      when "000010110111101" => color_data <= "100110000010";
      when "000010110111110" => color_data <= "011101100011";
      when "000010110111111" => color_data <= "010001000010";
      when "000010111000000" => color_data <= "000000000000";
      when "000010111000001" => color_data <= "000000000000";
      when "000010111000010" => color_data <= "000000000000";
      when "000010111000011" => color_data <= "000000000000";
      when "000010111000100" => color_data <= "000000000000";
      when "000010111000101" => color_data <= "000000000000";
      when "000010111000110" => color_data <= "000000000000";
      when "000010111000111" => color_data <= "000000000000";
      when "000010111001000" => color_data <= "000000000000";
      when "000010111001001" => color_data <= "000000000000";
      when "000010111001010" => color_data <= "000000000000";
      when "000010111001011" => color_data <= "000000000000";
      when "000010111001100" => color_data <= "000000000000";
      when "000010111001101" => color_data <= "000000000000";
      when "000010111001110" => color_data <= "000000000000";
      when "000010111001111" => color_data <= "000000000000";
      when "000010111010000" => color_data <= "000000000000";
      when "000010111010001" => color_data <= "000000000000";
      when "000010111010010" => color_data <= "000000000000";
      when "000010111010011" => color_data <= "000000000000";
      when "000010111010100" => color_data <= "000000000000";
      when "000010111010101" => color_data <= "000000000000";
      when "000010111010110" => color_data <= "000000000000";
      when "000010111010111" => color_data <= "000000000000";
      when "000010111011000" => color_data <= "000000000000";
      when "000010111011001" => color_data <= "000000000000";
      when "000010111011010" => color_data <= "000000000000";
      when "000010111011011" => color_data <= "000000000000";
      when "000010111011100" => color_data <= "000000000000";
      when "000010111011101" => color_data <= "000000000000";
      when "000010111011110" => color_data <= "000000000000";
      when "000010111011111" => color_data <= "000000000000";
      when "000010111100000" => color_data <= "000000000000";
      when "000010111100001" => color_data <= "000000000000";
      when "000010111100010" => color_data <= "000000000000";
      when "000010111100011" => color_data <= "000000000000";
      when "000011000000000" => color_data <= "000000000000";
      when "000011000000001" => color_data <= "000000000000";
      when "000011000000010" => color_data <= "000000000000";
      when "000011000000011" => color_data <= "000000000000";
      when "000011000000100" => color_data <= "000000000000";
      when "000011000000101" => color_data <= "000000000000";
      when "000011000000110" => color_data <= "000000000000";
      when "000011000000111" => color_data <= "000000000000";
      when "000011000001000" => color_data <= "000000000000";
      when "000011000001001" => color_data <= "000000000000";
      when "000011000001010" => color_data <= "000000000000";
      when "000011000001011" => color_data <= "000000000000";
      when "000011000001100" => color_data <= "000000000000";
      when "000011000001101" => color_data <= "000000000000";
      when "000011000001110" => color_data <= "000000000000";
      when "000011000001111" => color_data <= "000000000000";
      when "000011000010000" => color_data <= "000000000000";
      when "000011000010001" => color_data <= "000000000000";
      when "000011000010010" => color_data <= "000000000000";
      when "000011000010011" => color_data <= "000000000000";
      when "000011000010100" => color_data <= "000000000000";
      when "000011000010101" => color_data <= "000000000000";
      when "000011000010110" => color_data <= "000000000000";
      when "000011000010111" => color_data <= "000000000000";
      when "000011000011000" => color_data <= "000000000000";
      when "000011000011001" => color_data <= "000000000000";
      when "000011000011010" => color_data <= "000000000000";
      when "000011000011011" => color_data <= "000000000000";
      when "000011000011100" => color_data <= "000000000000";
      when "000011000011101" => color_data <= "000000000000";
      when "000011000011110" => color_data <= "000000000000";
      when "000011000011111" => color_data <= "000000000000";
      when "000011000100000" => color_data <= "000000000000";
      when "000011000100001" => color_data <= "000000000000";
      when "000011000100010" => color_data <= "000000000000";
      when "000011000100011" => color_data <= "010001000010";
      when "000011000100100" => color_data <= "100001110010";
      when "000011000100101" => color_data <= "111111010100";
      when "000011000100110" => color_data <= "111111100110";
      when "000011000100111" => color_data <= "111111101000";
      when "000011000101000" => color_data <= "111111010011";
      when "000011000101001" => color_data <= "111111010000";
      when "000011000101010" => color_data <= "111111010000";
      when "000011000101011" => color_data <= "111111010000";
      when "000011000101100" => color_data <= "111111010000";
      when "000011000101101" => color_data <= "111111010000";
      when "000011000101110" => color_data <= "111111010000";
      when "000011000101111" => color_data <= "111111010000";
      when "000011000110000" => color_data <= "111111010000";
      when "000011000110001" => color_data <= "111111010000";
      when "000011000110010" => color_data <= "111111010010";
      when "000011000110011" => color_data <= "111111100110";
      when "000011000110100" => color_data <= "111111010010";
      when "000011000110101" => color_data <= "111111010000";
      when "000011000110110" => color_data <= "111111010000";
      when "000011000110111" => color_data <= "111111010000";
      when "000011000111000" => color_data <= "111111010000";
      when "000011000111001" => color_data <= "111111010000";
      when "000011000111010" => color_data <= "111111010000";
      when "000011000111011" => color_data <= "111111010000";
      when "000011000111100" => color_data <= "111111010000";
      when "000011000111101" => color_data <= "111111010011";
      when "000011000111110" => color_data <= "111111100110";
      when "000011000111111" => color_data <= "100110000010";
      when "000011001000000" => color_data <= "011101110011";
      when "000011001000001" => color_data <= "001100110010";
      when "000011001000010" => color_data <= "000000000000";
      when "000011001000011" => color_data <= "000000000000";
      when "000011001000100" => color_data <= "000000000000";
      when "000011001000101" => color_data <= "000000000000";
      when "000011001000110" => color_data <= "000000000000";
      when "000011001000111" => color_data <= "000000000000";
      when "000011001001000" => color_data <= "000000000000";
      when "000011001001001" => color_data <= "000000000000";
      when "000011001001010" => color_data <= "000000000000";
      when "000011001001011" => color_data <= "000000000000";
      when "000011001001100" => color_data <= "000000000000";
      when "000011001001101" => color_data <= "000000000000";
      when "000011001001110" => color_data <= "000000000000";
      when "000011001001111" => color_data <= "000000000000";
      when "000011001010000" => color_data <= "000000000000";
      when "000011001010001" => color_data <= "000000000000";
      when "000011001010010" => color_data <= "000000000000";
      when "000011001010011" => color_data <= "000000000000";
      when "000011001010100" => color_data <= "000000000000";
      when "000011001010101" => color_data <= "000000000000";
      when "000011001010110" => color_data <= "000000000000";
      when "000011001010111" => color_data <= "000000000000";
      when "000011001011000" => color_data <= "000000000000";
      when "000011001011001" => color_data <= "000000000000";
      when "000011001011010" => color_data <= "000000000000";
      when "000011001011011" => color_data <= "000000000000";
      when "000011001011100" => color_data <= "000000000000";
      when "000011001011101" => color_data <= "000000000000";
      when "000011001011110" => color_data <= "000000000000";
      when "000011001011111" => color_data <= "000000000000";
      when "000011001100000" => color_data <= "000000000000";
      when "000011001100001" => color_data <= "000000000000";
      when "000011001100010" => color_data <= "000000000000";
      when "000011001100011" => color_data <= "000000000000";
      when "000011010000000" => color_data <= "000000000000";
      when "000011010000001" => color_data <= "000000000000";
      when "000011010000010" => color_data <= "000000000000";
      when "000011010000011" => color_data <= "000000000000";
      when "000011010000100" => color_data <= "000000000000";
      when "000011010000101" => color_data <= "000000000000";
      when "000011010000110" => color_data <= "000000000000";
      when "000011010000111" => color_data <= "000000000000";
      when "000011010001000" => color_data <= "000000000000";
      when "000011010001001" => color_data <= "000000000000";
      when "000011010001010" => color_data <= "000000000000";
      when "000011010001011" => color_data <= "000000000000";
      when "000011010001100" => color_data <= "000000000000";
      when "000011010001101" => color_data <= "000000000000";
      when "000011010001110" => color_data <= "000000000000";
      when "000011010001111" => color_data <= "000000000000";
      when "000011010010000" => color_data <= "000000000000";
      when "000011010010001" => color_data <= "000000000000";
      when "000011010010010" => color_data <= "000000000000";
      when "000011010010011" => color_data <= "000000000000";
      when "000011010010100" => color_data <= "000000000000";
      when "000011010010101" => color_data <= "000000000000";
      when "000011010010110" => color_data <= "000000000000";
      when "000011010010111" => color_data <= "000000000000";
      when "000011010011000" => color_data <= "000000000000";
      when "000011010011001" => color_data <= "000000000000";
      when "000011010011010" => color_data <= "000000000000";
      when "000011010011011" => color_data <= "000000000000";
      when "000011010011100" => color_data <= "000000000000";
      when "000011010011101" => color_data <= "000000000000";
      when "000011010011110" => color_data <= "000000000000";
      when "000011010011111" => color_data <= "000000000000";
      when "000011010100000" => color_data <= "000000000000";
      when "000011010100001" => color_data <= "001000100001";
      when "000011010100010" => color_data <= "100001110010";
      when "000011010100011" => color_data <= "100110000010";
      when "000011010100100" => color_data <= "111111100110";
      when "000011010100101" => color_data <= "111111101000";
      when "000011010100110" => color_data <= "111111100110";
      when "000011010100111" => color_data <= "111111010101";
      when "000011010101000" => color_data <= "111111010000";
      when "000011010101001" => color_data <= "111111000000";
      when "000011010101010" => color_data <= "111111010000";
      when "000011010101011" => color_data <= "111111010000";
      when "000011010101100" => color_data <= "111111010000";
      when "000011010101101" => color_data <= "111111010000";
      when "000011010101110" => color_data <= "111111010000";
      when "000011010101111" => color_data <= "111111010000";
      when "000011010110000" => color_data <= "111111010000";
      when "000011010110001" => color_data <= "111111010001";
      when "000011010110010" => color_data <= "111111010000";
      when "000011010110011" => color_data <= "111111010000";
      when "000011010110100" => color_data <= "111111010000";
      when "000011010110101" => color_data <= "111111010001";
      when "000011010110110" => color_data <= "111111010000";
      when "000011010110111" => color_data <= "111111010000";
      when "000011010111000" => color_data <= "111111010000";
      when "000011010111001" => color_data <= "111111010000";
      when "000011010111010" => color_data <= "111111010000";
      when "000011010111011" => color_data <= "111111010000";
      when "000011010111100" => color_data <= "111111010000";
      when "000011010111101" => color_data <= "111111010000";
      when "000011010111110" => color_data <= "111111100110";
      when "000011010111111" => color_data <= "111111101000";
      when "000011011000000" => color_data <= "111111100110";
      when "000011011000001" => color_data <= "100110000010";
      when "000011011000010" => color_data <= "011101110011";
      when "000011011000011" => color_data <= "000000000000";
      when "000011011000100" => color_data <= "000000000000";
      when "000011011000101" => color_data <= "000000000000";
      when "000011011000110" => color_data <= "000000000000";
      when "000011011000111" => color_data <= "000000000000";
      when "000011011001000" => color_data <= "000000000000";
      when "000011011001001" => color_data <= "000000000000";
      when "000011011001010" => color_data <= "000000000000";
      when "000011011001011" => color_data <= "000000000000";
      when "000011011001100" => color_data <= "000000000000";
      when "000011011001101" => color_data <= "000000000000";
      when "000011011001110" => color_data <= "000000000000";
      when "000011011001111" => color_data <= "000000000000";
      when "000011011010000" => color_data <= "000000000000";
      when "000011011010001" => color_data <= "000000000000";
      when "000011011010010" => color_data <= "000000000000";
      when "000011011010011" => color_data <= "000000000000";
      when "000011011010100" => color_data <= "000000000000";
      when "000011011010101" => color_data <= "000000000000";
      when "000011011010110" => color_data <= "000000000000";
      when "000011011010111" => color_data <= "000000000000";
      when "000011011011000" => color_data <= "000000000000";
      when "000011011011001" => color_data <= "000000000000";
      when "000011011011010" => color_data <= "000000000000";
      when "000011011011011" => color_data <= "000000000000";
      when "000011011011100" => color_data <= "000000000000";
      when "000011011011101" => color_data <= "000000000000";
      when "000011011011110" => color_data <= "000000000000";
      when "000011011011111" => color_data <= "000000000000";
      when "000011011100000" => color_data <= "000000000000";
      when "000011011100001" => color_data <= "000000000000";
      when "000011011100010" => color_data <= "000000000000";
      when "000011011100011" => color_data <= "000000000000";
      when "000011100000000" => color_data <= "000000000000";
      when "000011100000001" => color_data <= "000000000000";
      when "000011100000010" => color_data <= "000000000000";
      when "000011100000011" => color_data <= "000000000000";
      when "000011100000100" => color_data <= "000000000000";
      when "000011100000101" => color_data <= "000000000000";
      when "000011100000110" => color_data <= "000000000000";
      when "000011100000111" => color_data <= "000000000000";
      when "000011100001000" => color_data <= "000000000000";
      when "000011100001001" => color_data <= "000000000000";
      when "000011100001010" => color_data <= "000000000000";
      when "000011100001011" => color_data <= "000000000000";
      when "000011100001100" => color_data <= "000000000000";
      when "000011100001101" => color_data <= "000000000000";
      when "000011100001110" => color_data <= "000000000000";
      when "000011100001111" => color_data <= "000000000000";
      when "000011100010000" => color_data <= "000000000000";
      when "000011100010001" => color_data <= "000000000000";
      when "000011100010010" => color_data <= "000000000000";
      when "000011100010011" => color_data <= "000000000000";
      when "000011100010100" => color_data <= "000000000000";
      when "000011100010101" => color_data <= "000000000000";
      when "000011100010110" => color_data <= "000000000000";
      when "000011100010111" => color_data <= "000000000000";
      when "000011100011000" => color_data <= "000000000000";
      when "000011100011001" => color_data <= "000000000000";
      when "000011100011010" => color_data <= "000000000000";
      when "000011100011011" => color_data <= "000000000000";
      when "000011100011100" => color_data <= "000000000000";
      when "000011100011101" => color_data <= "000000000000";
      when "000011100011110" => color_data <= "000000000000";
      when "000011100011111" => color_data <= "000000000000";
      when "000011100100000" => color_data <= "010101010011";
      when "000011100100001" => color_data <= "100110000010";
      when "000011100100010" => color_data <= "111111100101";
      when "000011100100011" => color_data <= "111111101000";
      when "000011100100100" => color_data <= "111111100111";
      when "000011100100101" => color_data <= "111111010101";
      when "000011100100110" => color_data <= "111111100101";
      when "000011100100111" => color_data <= "111111111010";
      when "000011100101000" => color_data <= "111111111010";
      when "000011100101001" => color_data <= "111111010100";
      when "000011100101010" => color_data <= "111111000000";
      when "000011100101011" => color_data <= "111111000000";
      when "000011100101100" => color_data <= "111111010000";
      when "000011100101101" => color_data <= "111111010000";
      when "000011100101110" => color_data <= "111111010000";
      when "000011100101111" => color_data <= "111111010000";
      when "000011100110000" => color_data <= "111111010000";
      when "000011100110001" => color_data <= "111111010000";
      when "000011100110010" => color_data <= "111111010000";
      when "000011100110011" => color_data <= "111111010000";
      when "000011100110100" => color_data <= "111111010000";
      when "000011100110101" => color_data <= "111111010000";
      when "000011100110110" => color_data <= "111111010000";
      when "000011100110111" => color_data <= "111111010000";
      when "000011100111000" => color_data <= "111111010000";
      when "000011100111001" => color_data <= "111111010000";
      when "000011100111010" => color_data <= "111111010000";
      when "000011100111011" => color_data <= "111111010000";
      when "000011100111100" => color_data <= "111111010000";
      when "000011100111101" => color_data <= "111111000000";
      when "000011100111110" => color_data <= "111111010010";
      when "000011100111111" => color_data <= "111111100111";
      when "000011101000000" => color_data <= "111111100111";
      when "000011101000001" => color_data <= "111111100111";
      when "000011101000010" => color_data <= "111111010101";
      when "000011101000011" => color_data <= "100110000010";
      when "000011101000100" => color_data <= "001100110010";
      when "000011101000101" => color_data <= "000000000000";
      when "000011101000110" => color_data <= "000000000000";
      when "000011101000111" => color_data <= "000000000000";
      when "000011101001000" => color_data <= "000000000000";
      when "000011101001001" => color_data <= "000000000000";
      when "000011101001010" => color_data <= "000000000000";
      when "000011101001011" => color_data <= "000000000000";
      when "000011101001100" => color_data <= "000000000000";
      when "000011101001101" => color_data <= "000000000000";
      when "000011101001110" => color_data <= "000000000000";
      when "000011101001111" => color_data <= "000000000000";
      when "000011101010000" => color_data <= "000000000000";
      when "000011101010001" => color_data <= "000000000000";
      when "000011101010010" => color_data <= "000000000000";
      when "000011101010011" => color_data <= "000000000000";
      when "000011101010100" => color_data <= "000000000000";
      when "000011101010101" => color_data <= "000000000000";
      when "000011101010110" => color_data <= "000000000000";
      when "000011101010111" => color_data <= "000000000000";
      when "000011101011000" => color_data <= "000000000000";
      when "000011101011001" => color_data <= "000000000000";
      when "000011101011010" => color_data <= "000000000000";
      when "000011101011011" => color_data <= "000000000000";
      when "000011101011100" => color_data <= "000000000000";
      when "000011101011101" => color_data <= "000000000000";
      when "000011101011110" => color_data <= "000000000000";
      when "000011101011111" => color_data <= "000000000000";
      when "000011101100000" => color_data <= "000000000000";
      when "000011101100001" => color_data <= "000000000000";
      when "000011101100010" => color_data <= "000000000000";
      when "000011101100011" => color_data <= "000000000000";
      when "000011110000000" => color_data <= "000000000000";
      when "000011110000001" => color_data <= "000000000000";
      when "000011110000010" => color_data <= "000000000000";
      when "000011110000011" => color_data <= "000000000000";
      when "000011110000100" => color_data <= "000000000000";
      when "000011110000101" => color_data <= "000000000000";
      when "000011110000110" => color_data <= "000000000000";
      when "000011110000111" => color_data <= "000000000000";
      when "000011110001000" => color_data <= "000000000000";
      when "000011110001001" => color_data <= "000000000000";
      when "000011110001010" => color_data <= "000000000000";
      when "000011110001011" => color_data <= "000000000000";
      when "000011110001100" => color_data <= "000000000000";
      when "000011110001101" => color_data <= "000000000000";
      when "000011110001110" => color_data <= "000000000000";
      when "000011110001111" => color_data <= "000000000000";
      when "000011110010000" => color_data <= "000000000000";
      when "000011110010001" => color_data <= "000000000000";
      when "000011110010010" => color_data <= "000000000000";
      when "000011110010011" => color_data <= "000000000000";
      when "000011110010100" => color_data <= "000000000000";
      when "000011110010101" => color_data <= "000000000000";
      when "000011110010110" => color_data <= "000000000000";
      when "000011110010111" => color_data <= "000000000000";
      when "000011110011000" => color_data <= "000000000000";
      when "000011110011001" => color_data <= "000000000000";
      when "000011110011010" => color_data <= "000000000000";
      when "000011110011011" => color_data <= "000000000000";
      when "000011110011100" => color_data <= "000000000000";
      when "000011110011101" => color_data <= "000000000000";
      when "000011110011110" => color_data <= "000000000000";
      when "000011110011111" => color_data <= "011101110011";
      when "000011110100000" => color_data <= "100110000010";
      when "000011110100001" => color_data <= "111111100111";
      when "000011110100010" => color_data <= "111111100111";
      when "000011110100011" => color_data <= "111111100110";
      when "000011110100100" => color_data <= "111111010100";
      when "000011110100101" => color_data <= "111111100111";
      when "000011110100110" => color_data <= "111111111100";
      when "000011110100111" => color_data <= "111111111110";
      when "000011110101000" => color_data <= "111111111111";
      when "000011110101001" => color_data <= "111111111110";
      when "000011110101010" => color_data <= "111111111011";
      when "000011110101011" => color_data <= "111111100101";
      when "000011110101100" => color_data <= "111111010000";
      when "000011110101101" => color_data <= "111111000000";
      when "000011110101110" => color_data <= "111111010000";
      when "000011110101111" => color_data <= "111111010000";
      when "000011110110000" => color_data <= "111111010000";
      when "000011110110001" => color_data <= "111111010000";
      when "000011110110010" => color_data <= "111111010000";
      when "000011110110011" => color_data <= "111111010000";
      when "000011110110100" => color_data <= "111111010000";
      when "000011110110101" => color_data <= "111111010000";
      when "000011110110110" => color_data <= "111111010000";
      when "000011110110111" => color_data <= "111111010000";
      when "000011110111000" => color_data <= "111111010000";
      when "000011110111001" => color_data <= "111111010000";
      when "000011110111010" => color_data <= "111111010000";
      when "000011110111011" => color_data <= "111111010000";
      when "000011110111100" => color_data <= "111111010010";
      when "000011110111101" => color_data <= "111111010011";
      when "000011110111110" => color_data <= "111111100101";
      when "000011110111111" => color_data <= "111111100100";
      when "000011111000000" => color_data <= "111111100101";
      when "000011111000001" => color_data <= "111111100111";
      when "000011111000010" => color_data <= "111111101000";
      when "000011111000011" => color_data <= "111111100110";
      when "000011111000100" => color_data <= "100110000010";
      when "000011111000101" => color_data <= "010101010011";
      when "000011111000110" => color_data <= "000000000000";
      when "000011111000111" => color_data <= "000000000000";
      when "000011111001000" => color_data <= "000000000000";
      when "000011111001001" => color_data <= "000000000000";
      when "000011111001010" => color_data <= "000000000000";
      when "000011111001011" => color_data <= "000000000000";
      when "000011111001100" => color_data <= "000000000000";
      when "000011111001101" => color_data <= "000000000000";
      when "000011111001110" => color_data <= "000000000000";
      when "000011111001111" => color_data <= "000000000000";
      when "000011111010000" => color_data <= "000000000000";
      when "000011111010001" => color_data <= "000000000000";
      when "000011111010010" => color_data <= "000000000000";
      when "000011111010011" => color_data <= "000000000000";
      when "000011111010100" => color_data <= "000000000000";
      when "000011111010101" => color_data <= "000000000000";
      when "000011111010110" => color_data <= "000000000000";
      when "000011111010111" => color_data <= "000000000000";
      when "000011111011000" => color_data <= "000000000000";
      when "000011111011001" => color_data <= "000000000000";
      when "000011111011010" => color_data <= "000000000000";
      when "000011111011011" => color_data <= "000000000000";
      when "000011111011100" => color_data <= "000000000000";
      when "000011111011101" => color_data <= "000000000000";
      when "000011111011110" => color_data <= "000000000000";
      when "000011111011111" => color_data <= "000000000000";
      when "000011111100000" => color_data <= "000000000000";
      when "000011111100001" => color_data <= "000000000000";
      when "000011111100010" => color_data <= "000000000000";
      when "000011111100011" => color_data <= "000000000000";
      when "000100000000000" => color_data <= "000000000000";
      when "000100000000001" => color_data <= "000000000000";
      when "000100000000010" => color_data <= "000000000000";
      when "000100000000011" => color_data <= "000000000000";
      when "000100000000100" => color_data <= "000000000000";
      when "000100000000101" => color_data <= "000000000000";
      when "000100000000110" => color_data <= "000000000000";
      when "000100000000111" => color_data <= "000000000000";
      when "000100000001000" => color_data <= "000000000000";
      when "000100000001001" => color_data <= "000000000000";
      when "000100000001010" => color_data <= "000000000000";
      when "000100000001011" => color_data <= "000000000000";
      when "000100000001100" => color_data <= "000000000000";
      when "000100000001101" => color_data <= "000000000000";
      when "000100000001110" => color_data <= "000000000000";
      when "000100000001111" => color_data <= "000000000000";
      when "000100000010000" => color_data <= "000000000000";
      when "000100000010001" => color_data <= "000000000000";
      when "000100000010010" => color_data <= "000000000000";
      when "000100000010011" => color_data <= "000000000000";
      when "000100000010100" => color_data <= "000000000000";
      when "000100000010101" => color_data <= "000000000000";
      when "000100000010110" => color_data <= "000000000000";
      when "000100000010111" => color_data <= "000000000000";
      when "000100000011000" => color_data <= "000000000000";
      when "000100000011001" => color_data <= "000000000000";
      when "000100000011010" => color_data <= "000000000000";
      when "000100000011011" => color_data <= "000000000000";
      when "000100000011100" => color_data <= "000000000000";
      when "000100000011101" => color_data <= "000000000000";
      when "000100000011110" => color_data <= "100010000010";
      when "000100000011111" => color_data <= "100001110010";
      when "000100000100000" => color_data <= "111111100111";
      when "000100000100001" => color_data <= "111111100111";
      when "000100000100010" => color_data <= "111111100101";
      when "000100000100011" => color_data <= "111111100101";
      when "000100000100100" => color_data <= "111111111010";
      when "000100000100101" => color_data <= "111111111110";
      when "000100000100110" => color_data <= "111111111101";
      when "000100000100111" => color_data <= "111111111101";
      when "000100000101000" => color_data <= "111111111100";
      when "000100000101001" => color_data <= "111111111101";
      when "000100000101010" => color_data <= "111111111110";
      when "000100000101011" => color_data <= "111111111111";
      when "000100000101100" => color_data <= "111111111011";
      when "000100000101101" => color_data <= "111111100110";
      when "000100000101110" => color_data <= "111111010001";
      when "000100000101111" => color_data <= "111111000000";
      when "000100000110000" => color_data <= "111111010000";
      when "000100000110001" => color_data <= "111111010000";
      when "000100000110010" => color_data <= "111111010000";
      when "000100000110011" => color_data <= "111111010000";
      when "000100000110100" => color_data <= "111111010001";
      when "000100000110101" => color_data <= "111111010000";
      when "000100000110110" => color_data <= "111111010000";
      when "000100000110111" => color_data <= "111111010000";
      when "000100000111000" => color_data <= "111111010000";
      when "000100000111001" => color_data <= "111111010010";
      when "000100000111010" => color_data <= "111111010100";
      when "000100000111011" => color_data <= "111111100110";
      when "000100000111100" => color_data <= "111111100111";
      when "000100000111101" => color_data <= "111111101000";
      when "000100000111110" => color_data <= "111111101000";
      when "000100000111111" => color_data <= "111111100110";
      when "000100001000000" => color_data <= "111111010100";
      when "000100001000001" => color_data <= "111111010100";
      when "000100001000010" => color_data <= "111111100110";
      when "000100001000011" => color_data <= "111111100111";
      when "000100001000100" => color_data <= "111111100111";
      when "000100001000101" => color_data <= "100110000010";
      when "000100001000110" => color_data <= "011101100011";
      when "000100001000111" => color_data <= "000000000000";
      when "000100001001000" => color_data <= "000000000000";
      when "000100001001001" => color_data <= "000000000000";
      when "000100001001010" => color_data <= "000000000000";
      when "000100001001011" => color_data <= "000000000000";
      when "000100001001100" => color_data <= "000000000000";
      when "000100001001101" => color_data <= "000000000000";
      when "000100001001110" => color_data <= "000000000000";
      when "000100001001111" => color_data <= "000000000000";
      when "000100001010000" => color_data <= "000000000000";
      when "000100001010001" => color_data <= "000000000000";
      when "000100001010010" => color_data <= "000000000000";
      when "000100001010011" => color_data <= "000000000000";
      when "000100001010100" => color_data <= "000000000000";
      when "000100001010101" => color_data <= "000000000000";
      when "000100001010110" => color_data <= "000000000000";
      when "000100001010111" => color_data <= "000000000000";
      when "000100001011000" => color_data <= "000000000000";
      when "000100001011001" => color_data <= "000000000000";
      when "000100001011010" => color_data <= "000000000000";
      when "000100001011011" => color_data <= "000000000000";
      when "000100001011100" => color_data <= "000000000000";
      when "000100001011101" => color_data <= "000000000000";
      when "000100001011110" => color_data <= "000000000000";
      when "000100001011111" => color_data <= "000000000000";
      when "000100001100000" => color_data <= "000000000000";
      when "000100001100001" => color_data <= "000000000000";
      when "000100001100010" => color_data <= "000000000000";
      when "000100001100011" => color_data <= "000000000000";
      when "000100010000000" => color_data <= "000000000000";
      when "000100010000001" => color_data <= "000000000000";
      when "000100010000010" => color_data <= "000000000000";
      when "000100010000011" => color_data <= "000000000000";
      when "000100010000100" => color_data <= "000000000000";
      when "000100010000101" => color_data <= "000000000000";
      when "000100010000110" => color_data <= "000000000000";
      when "000100010000111" => color_data <= "000000000000";
      when "000100010001000" => color_data <= "000000000000";
      when "000100010001001" => color_data <= "000000000000";
      when "000100010001010" => color_data <= "000000000000";
      when "000100010001011" => color_data <= "000000000000";
      when "000100010001100" => color_data <= "000000000000";
      when "000100010001101" => color_data <= "000000000000";
      when "000100010001110" => color_data <= "000000000000";
      when "000100010001111" => color_data <= "000000000000";
      when "000100010010000" => color_data <= "000000000000";
      when "000100010010001" => color_data <= "000000000000";
      when "000100010010010" => color_data <= "000000000000";
      when "000100010010011" => color_data <= "000000000000";
      when "000100010010100" => color_data <= "000000000000";
      when "000100010010101" => color_data <= "000000000000";
      when "000100010010110" => color_data <= "000000000000";
      when "000100010010111" => color_data <= "000000000000";
      when "000100010011000" => color_data <= "000000000000";
      when "000100010011001" => color_data <= "000000000000";
      when "000100010011010" => color_data <= "000000000000";
      when "000100010011011" => color_data <= "000000000000";
      when "000100010011100" => color_data <= "000000000000";
      when "000100010011101" => color_data <= "100110000010";
      when "000100010011110" => color_data <= "111111100101";
      when "000100010011111" => color_data <= "111111101000";
      when "000100010100000" => color_data <= "111111100110";
      when "000100010100001" => color_data <= "111111010100";
      when "000100010100010" => color_data <= "111111100111";
      when "000100010100011" => color_data <= "111111111101";
      when "000100010100100" => color_data <= "111111111110";
      when "000100010100101" => color_data <= "111111111101";
      when "000100010100110" => color_data <= "111111111100";
      when "000100010100111" => color_data <= "111111111101";
      when "000100010101000" => color_data <= "111111111101";
      when "000100010101001" => color_data <= "111111111101";
      when "000100010101010" => color_data <= "111111111100";
      when "000100010101011" => color_data <= "111111111101";
      when "000100010101100" => color_data <= "111111111110";
      when "000100010101101" => color_data <= "111111111111";
      when "000100010101110" => color_data <= "111111111100";
      when "000100010101111" => color_data <= "111111100111";
      when "000100010110000" => color_data <= "111111010010";
      when "000100010110001" => color_data <= "111111000000";
      when "000100010110010" => color_data <= "111111010000";
      when "000100010110011" => color_data <= "111111010000";
      when "000100010110100" => color_data <= "111111010000";
      when "000100010110101" => color_data <= "111111010000";
      when "000100010110110" => color_data <= "111111010001";
      when "000100010110111" => color_data <= "111111010100";
      when "000100010111000" => color_data <= "111111100110";
      when "000100010111001" => color_data <= "111111100111";
      when "000100010111010" => color_data <= "111111101000";
      when "000100010111011" => color_data <= "111111100111";
      when "000100010111100" => color_data <= "111111100111";
      when "000100010111101" => color_data <= "111111100111";
      when "000100010111110" => color_data <= "111111100110";
      when "000100010111111" => color_data <= "111111100111";
      when "000100011000000" => color_data <= "111111100111";
      when "000100011000001" => color_data <= "111111100110";
      when "000100011000010" => color_data <= "111111010100";
      when "000100011000011" => color_data <= "111111010101";
      when "000100011000100" => color_data <= "111111100111";
      when "000100011000101" => color_data <= "111111101000";
      when "000100011000110" => color_data <= "100110000010";
      when "000100011000111" => color_data <= "011101110011";
      when "000100011001000" => color_data <= "000000000000";
      when "000100011001001" => color_data <= "000000000000";
      when "000100011001010" => color_data <= "000000000000";
      when "000100011001011" => color_data <= "000000000000";
      when "000100011001100" => color_data <= "000000000000";
      when "000100011001101" => color_data <= "000000000000";
      when "000100011001110" => color_data <= "000000000000";
      when "000100011001111" => color_data <= "000000000000";
      when "000100011010000" => color_data <= "000000000000";
      when "000100011010001" => color_data <= "000000000000";
      when "000100011010010" => color_data <= "000000000000";
      when "000100011010011" => color_data <= "000000000000";
      when "000100011010100" => color_data <= "000000000000";
      when "000100011010101" => color_data <= "000000000000";
      when "000100011010110" => color_data <= "000000000000";
      when "000100011010111" => color_data <= "000000000000";
      when "000100011011000" => color_data <= "000000000000";
      when "000100011011001" => color_data <= "000000000000";
      when "000100011011010" => color_data <= "000000000000";
      when "000100011011011" => color_data <= "000000000000";
      when "000100011011100" => color_data <= "000000000000";
      when "000100011011101" => color_data <= "000000000000";
      when "000100011011110" => color_data <= "000000000000";
      when "000100011011111" => color_data <= "000000000000";
      when "000100011100000" => color_data <= "000000000000";
      when "000100011100001" => color_data <= "000000000000";
      when "000100011100010" => color_data <= "000000000000";
      when "000100011100011" => color_data <= "000000000000";
      when "000100100000000" => color_data <= "000000000000";
      when "000100100000001" => color_data <= "000000000000";
      when "000100100000010" => color_data <= "000000000000";
      when "000100100000011" => color_data <= "000000000000";
      when "000100100000100" => color_data <= "000000000000";
      when "000100100000101" => color_data <= "000000000000";
      when "000100100000110" => color_data <= "000000000000";
      when "000100100000111" => color_data <= "000000000000";
      when "000100100001000" => color_data <= "000000000000";
      when "000100100001001" => color_data <= "000000000000";
      when "000100100001010" => color_data <= "000000000000";
      when "000100100001011" => color_data <= "000000000000";
      when "000100100001100" => color_data <= "000000000000";
      when "000100100001101" => color_data <= "000000000000";
      when "000100100001110" => color_data <= "000000000000";
      when "000100100001111" => color_data <= "000000000000";
      when "000100100010000" => color_data <= "000000000000";
      when "000100100010001" => color_data <= "000000000000";
      when "000100100010010" => color_data <= "000000000000";
      when "000100100010011" => color_data <= "000000000000";
      when "000100100010100" => color_data <= "000000000000";
      when "000100100010101" => color_data <= "000000000000";
      when "000100100010110" => color_data <= "000000000000";
      when "000100100010111" => color_data <= "000000000000";
      when "000100100011000" => color_data <= "000000000000";
      when "000100100011001" => color_data <= "000000000000";
      when "000100100011010" => color_data <= "000000000000";
      when "000100100011011" => color_data <= "000000000000";
      when "000100100011100" => color_data <= "100110000010";
      when "000100100011101" => color_data <= "111111100101";
      when "000100100011110" => color_data <= "111111101000";
      when "000100100011111" => color_data <= "111111100110";
      when "000100100100000" => color_data <= "111111010100";
      when "000100100100001" => color_data <= "111111101001";
      when "000100100100010" => color_data <= "111111111110";
      when "000100100100011" => color_data <= "111111111110";
      when "000100100100100" => color_data <= "111111111100";
      when "000100100100101" => color_data <= "111111111101";
      when "000100100100110" => color_data <= "111111111101";
      when "000100100100111" => color_data <= "111111111101";
      when "000100100101000" => color_data <= "111111111101";
      when "000100100101001" => color_data <= "111111111101";
      when "000100100101010" => color_data <= "111111111101";
      when "000100100101011" => color_data <= "111111111101";
      when "000100100101100" => color_data <= "111111111101";
      when "000100100101101" => color_data <= "111111111101";
      when "000100100101110" => color_data <= "111111111110";
      when "000100100101111" => color_data <= "111111111111";
      when "000100100110000" => color_data <= "111111111101";
      when "000100100110001" => color_data <= "111111101000";
      when "000100100110010" => color_data <= "111111010010";
      when "000100100110011" => color_data <= "111111010000";
      when "000100100110100" => color_data <= "111111010010";
      when "000100100110101" => color_data <= "111111010101";
      when "000100100110110" => color_data <= "111111100111";
      when "000100100110111" => color_data <= "111111101000";
      when "000100100111000" => color_data <= "111111100111";
      when "000100100111001" => color_data <= "111111100111";
      when "000100100111010" => color_data <= "111111100111";
      when "000100100111011" => color_data <= "111111100111";
      when "000100100111100" => color_data <= "111111100111";
      when "000100100111101" => color_data <= "111111100111";
      when "000100100111110" => color_data <= "111111100111";
      when "000100100111111" => color_data <= "111111100111";
      when "000100101000000" => color_data <= "111111100111";
      when "000100101000001" => color_data <= "111111100111";
      when "000100101000010" => color_data <= "111111100111";
      when "000100101000011" => color_data <= "111111100101";
      when "000100101000100" => color_data <= "111111010100";
      when "000100101000101" => color_data <= "111111100110";
      when "000100101000110" => color_data <= "111111101000";
      when "000100101000111" => color_data <= "100110000010";
      when "000100101001000" => color_data <= "011101100011";
      when "000100101001001" => color_data <= "000000000000";
      when "000100101001010" => color_data <= "000000000000";
      when "000100101001011" => color_data <= "000000000000";
      when "000100101001100" => color_data <= "000000000000";
      when "000100101001101" => color_data <= "000000000000";
      when "000100101001110" => color_data <= "000000000000";
      when "000100101001111" => color_data <= "000000000000";
      when "000100101010000" => color_data <= "000000000000";
      when "000100101010001" => color_data <= "000000000000";
      when "000100101010010" => color_data <= "000000000000";
      when "000100101010011" => color_data <= "000000000000";
      when "000100101010100" => color_data <= "000000000000";
      when "000100101010101" => color_data <= "000000000000";
      when "000100101010110" => color_data <= "000000000000";
      when "000100101010111" => color_data <= "000000000000";
      when "000100101011000" => color_data <= "000000000000";
      when "000100101011001" => color_data <= "000000000000";
      when "000100101011010" => color_data <= "000000000000";
      when "000100101011011" => color_data <= "000000000000";
      when "000100101011100" => color_data <= "000000000000";
      when "000100101011101" => color_data <= "000000000000";
      when "000100101011110" => color_data <= "000000000000";
      when "000100101011111" => color_data <= "000000000000";
      when "000100101100000" => color_data <= "000000000000";
      when "000100101100001" => color_data <= "000000000000";
      when "000100101100010" => color_data <= "000000000000";
      when "000100101100011" => color_data <= "000000000000";
      when "000100110000000" => color_data <= "000000000000";
      when "000100110000001" => color_data <= "000000000000";
      when "000100110000010" => color_data <= "000000000000";
      when "000100110000011" => color_data <= "000000000000";
      when "000100110000100" => color_data <= "000000000000";
      when "000100110000101" => color_data <= "000000000000";
      when "000100110000110" => color_data <= "000000000000";
      when "000100110000111" => color_data <= "000000000000";
      when "000100110001000" => color_data <= "000000000000";
      when "000100110001001" => color_data <= "000000000000";
      when "000100110001010" => color_data <= "000000000000";
      when "000100110001011" => color_data <= "000000000000";
      when "000100110001100" => color_data <= "000000000000";
      when "000100110001101" => color_data <= "000000000000";
      when "000100110001110" => color_data <= "000000000000";
      when "000100110001111" => color_data <= "000000000000";
      when "000100110010000" => color_data <= "000000000000";
      when "000100110010001" => color_data <= "000000000000";
      when "000100110010010" => color_data <= "000000000000";
      when "000100110010011" => color_data <= "000000000000";
      when "000100110010100" => color_data <= "000000000000";
      when "000100110010101" => color_data <= "000000000000";
      when "000100110010110" => color_data <= "000000000000";
      when "000100110010111" => color_data <= "000000000000";
      when "000100110011000" => color_data <= "000000000000";
      when "000100110011001" => color_data <= "000000000000";
      when "000100110011010" => color_data <= "000000000000";
      when "000100110011011" => color_data <= "100001110010";
      when "000100110011100" => color_data <= "111111100101";
      when "000100110011101" => color_data <= "111111101000";
      when "000100110011110" => color_data <= "111111100101";
      when "000100110011111" => color_data <= "111111010100";
      when "000100110100000" => color_data <= "111111111010";
      when "000100110100001" => color_data <= "111111111110";
      when "000100110100010" => color_data <= "111111111101";
      when "000100110100011" => color_data <= "111111111100";
      when "000100110100100" => color_data <= "111111111101";
      when "000100110100101" => color_data <= "111111111101";
      when "000100110100110" => color_data <= "111111111101";
      when "000100110100111" => color_data <= "111111111101";
      when "000100110101000" => color_data <= "111111111101";
      when "000100110101001" => color_data <= "111111111101";
      when "000100110101010" => color_data <= "111111111101";
      when "000100110101011" => color_data <= "111111111101";
      when "000100110101100" => color_data <= "111111111101";
      when "000100110101101" => color_data <= "111111111101";
      when "000100110101110" => color_data <= "111111111101";
      when "000100110101111" => color_data <= "111111111100";
      when "000100110110000" => color_data <= "111111111101";
      when "000100110110001" => color_data <= "111111111111";
      when "000100110110010" => color_data <= "111111101001";
      when "000100110110011" => color_data <= "111111010100";
      when "000100110110100" => color_data <= "111111100111";
      when "000100110110101" => color_data <= "111111101000";
      when "000100110110110" => color_data <= "111111100111";
      when "000100110110111" => color_data <= "111111100111";
      when "000100110111000" => color_data <= "111111100111";
      when "000100110111001" => color_data <= "111111100111";
      when "000100110111010" => color_data <= "111111100111";
      when "000100110111011" => color_data <= "111111100111";
      when "000100110111100" => color_data <= "111111100111";
      when "000100110111101" => color_data <= "111111100111";
      when "000100110111110" => color_data <= "111111100111";
      when "000100110111111" => color_data <= "111111100111";
      when "000100111000000" => color_data <= "111111100111";
      when "000100111000001" => color_data <= "111111100111";
      when "000100111000010" => color_data <= "111111100111";
      when "000100111000011" => color_data <= "111111100111";
      when "000100111000100" => color_data <= "111111100110";
      when "000100111000101" => color_data <= "111111010100";
      when "000100111000110" => color_data <= "111111100110";
      when "000100111000111" => color_data <= "111111101000";
      when "000100111001000" => color_data <= "100110000010";
      when "000100111001001" => color_data <= "011001100011";
      when "000100111001010" => color_data <= "000000000000";
      when "000100111001011" => color_data <= "000000000000";
      when "000100111001100" => color_data <= "000000000000";
      when "000100111001101" => color_data <= "000000000000";
      when "000100111001110" => color_data <= "000000000000";
      when "000100111001111" => color_data <= "000000000000";
      when "000100111010000" => color_data <= "000000000000";
      when "000100111010001" => color_data <= "000000000000";
      when "000100111010010" => color_data <= "000000000000";
      when "000100111010011" => color_data <= "000000000000";
      when "000100111010100" => color_data <= "000000000000";
      when "000100111010101" => color_data <= "000000000000";
      when "000100111010110" => color_data <= "000000000000";
      when "000100111010111" => color_data <= "000000000000";
      when "000100111011000" => color_data <= "000000000000";
      when "000100111011001" => color_data <= "000000000000";
      when "000100111011010" => color_data <= "000000000000";
      when "000100111011011" => color_data <= "000000000000";
      when "000100111011100" => color_data <= "000000000000";
      when "000100111011101" => color_data <= "000000000000";
      when "000100111011110" => color_data <= "000000000000";
      when "000100111011111" => color_data <= "000000000000";
      when "000100111100000" => color_data <= "000000000000";
      when "000100111100001" => color_data <= "000000000000";
      when "000100111100010" => color_data <= "000000000000";
      when "000100111100011" => color_data <= "000000000000";
      when "000101000000000" => color_data <= "000000000000";
      when "000101000000001" => color_data <= "000000000000";
      when "000101000000010" => color_data <= "000000000000";
      when "000101000000011" => color_data <= "000000000000";
      when "000101000000100" => color_data <= "000000000000";
      when "000101000000101" => color_data <= "000000000000";
      when "000101000000110" => color_data <= "000000000000";
      when "000101000000111" => color_data <= "000000000000";
      when "000101000001000" => color_data <= "000000000000";
      when "000101000001001" => color_data <= "000000000000";
      when "000101000001010" => color_data <= "000000000000";
      when "000101000001011" => color_data <= "000000000000";
      when "000101000001100" => color_data <= "000000000000";
      when "000101000001101" => color_data <= "000000000000";
      when "000101000001110" => color_data <= "000000000000";
      when "000101000001111" => color_data <= "000000000000";
      when "000101000010000" => color_data <= "000000000000";
      when "000101000010001" => color_data <= "000000000000";
      when "000101000010010" => color_data <= "000000000000";
      when "000101000010011" => color_data <= "000000000000";
      when "000101000010100" => color_data <= "000000000000";
      when "000101000010101" => color_data <= "000000000000";
      when "000101000010110" => color_data <= "000000000000";
      when "000101000010111" => color_data <= "000000000000";
      when "000101000011000" => color_data <= "000000000000";
      when "000101000011001" => color_data <= "000000000000";
      when "000101000011010" => color_data <= "011001100011";
      when "000101000011011" => color_data <= "100001110011";
      when "000101000011100" => color_data <= "111111101001";
      when "000101000011101" => color_data <= "111111010101";
      when "000101000011110" => color_data <= "111111100101";
      when "000101000011111" => color_data <= "111111111100";
      when "000101000100000" => color_data <= "111111111110";
      when "000101000100001" => color_data <= "111111111101";
      when "000101000100010" => color_data <= "111111111101";
      when "000101000100011" => color_data <= "111111111101";
      when "000101000100100" => color_data <= "111111111101";
      when "000101000100101" => color_data <= "111111111101";
      when "000101000100110" => color_data <= "111111111101";
      when "000101000100111" => color_data <= "111111111101";
      when "000101000101000" => color_data <= "111111111101";
      when "000101000101001" => color_data <= "111111111101";
      when "000101000101010" => color_data <= "111111111101";
      when "000101000101011" => color_data <= "111111111101";
      when "000101000101100" => color_data <= "111111111101";
      when "000101000101101" => color_data <= "111111111101";
      when "000101000101110" => color_data <= "111111111101";
      when "000101000101111" => color_data <= "111111111101";
      when "000101000110000" => color_data <= "111111111101";
      when "000101000110001" => color_data <= "111111111110";
      when "000101000110010" => color_data <= "111111101001";
      when "000101000110011" => color_data <= "111111100101";
      when "000101000110100" => color_data <= "111111100111";
      when "000101000110101" => color_data <= "111111100111";
      when "000101000110110" => color_data <= "111111100111";
      when "000101000110111" => color_data <= "111111100111";
      when "000101000111000" => color_data <= "111111100111";
      when "000101000111001" => color_data <= "111111100111";
      when "000101000111010" => color_data <= "111111100111";
      when "000101000111011" => color_data <= "111111100111";
      when "000101000111100" => color_data <= "111111100111";
      when "000101000111101" => color_data <= "111111100111";
      when "000101000111110" => color_data <= "111111100111";
      when "000101000111111" => color_data <= "111111100111";
      when "000101001000000" => color_data <= "111111100111";
      when "000101001000001" => color_data <= "111111100111";
      when "000101001000010" => color_data <= "111111100111";
      when "000101001000011" => color_data <= "111111100111";
      when "000101001000100" => color_data <= "111111100111";
      when "000101001000101" => color_data <= "111111100110";
      when "000101001000110" => color_data <= "111111010100";
      when "000101001000111" => color_data <= "111111100101";
      when "000101001001000" => color_data <= "111111101000";
      when "000101001001001" => color_data <= "100110000010";
      when "000101001001010" => color_data <= "010001000010";
      when "000101001001011" => color_data <= "000000000000";
      when "000101001001100" => color_data <= "000000000000";
      when "000101001001101" => color_data <= "000000000000";
      when "000101001001110" => color_data <= "000000000000";
      when "000101001001111" => color_data <= "000000000000";
      when "000101001010000" => color_data <= "000000000000";
      when "000101001010001" => color_data <= "000000000000";
      when "000101001010010" => color_data <= "000000000000";
      when "000101001010011" => color_data <= "000000000000";
      when "000101001010100" => color_data <= "000000000000";
      when "000101001010101" => color_data <= "000000000000";
      when "000101001010110" => color_data <= "000000000000";
      when "000101001010111" => color_data <= "000000000000";
      when "000101001011000" => color_data <= "000000000000";
      when "000101001011001" => color_data <= "000000000000";
      when "000101001011010" => color_data <= "000000000000";
      when "000101001011011" => color_data <= "000000000000";
      when "000101001011100" => color_data <= "000000000000";
      when "000101001011101" => color_data <= "000000000000";
      when "000101001011110" => color_data <= "000000000000";
      when "000101001011111" => color_data <= "000000000000";
      when "000101001100000" => color_data <= "000000000000";
      when "000101001100001" => color_data <= "000000000000";
      when "000101001100010" => color_data <= "000000000000";
      when "000101001100011" => color_data <= "000000000000";
      when "000101010000000" => color_data <= "000000000000";
      when "000101010000001" => color_data <= "000000000000";
      when "000101010000010" => color_data <= "000000000000";
      when "000101010000011" => color_data <= "000000000000";
      when "000101010000100" => color_data <= "000000000000";
      when "000101010000101" => color_data <= "000000000000";
      when "000101010000110" => color_data <= "000000000000";
      when "000101010000111" => color_data <= "000000000000";
      when "000101010001000" => color_data <= "000000000000";
      when "000101010001001" => color_data <= "000000000000";
      when "000101010001010" => color_data <= "000000000000";
      when "000101010001011" => color_data <= "000000000000";
      when "000101010001100" => color_data <= "000000000000";
      when "000101010001101" => color_data <= "000000000000";
      when "000101010001110" => color_data <= "000000000000";
      when "000101010001111" => color_data <= "000000000000";
      when "000101010010000" => color_data <= "000000000000";
      when "000101010010001" => color_data <= "000000000000";
      when "000101010010010" => color_data <= "000000000000";
      when "000101010010011" => color_data <= "000000000000";
      when "000101010010100" => color_data <= "000000000000";
      when "000101010010101" => color_data <= "000000000000";
      when "000101010010110" => color_data <= "000000000000";
      when "000101010010111" => color_data <= "000000000000";
      when "000101010011000" => color_data <= "000000000000";
      when "000101010011001" => color_data <= "010101000010";
      when "000101010011010" => color_data <= "110110110000";
      when "000101010011011" => color_data <= "111111010100";
      when "000101010011100" => color_data <= "111111010011";
      when "000101010011101" => color_data <= "111111100110";
      when "000101010011110" => color_data <= "111111111101";
      when "000101010011111" => color_data <= "111111111110";
      when "000101010100000" => color_data <= "111111111101";
      when "000101010100001" => color_data <= "111111111101";
      when "000101010100010" => color_data <= "111111111101";
      when "000101010100011" => color_data <= "111111111101";
      when "000101010100100" => color_data <= "111111111101";
      when "000101010100101" => color_data <= "111111111101";
      when "000101010100110" => color_data <= "111111111101";
      when "000101010100111" => color_data <= "111111111101";
      when "000101010101000" => color_data <= "111111111101";
      when "000101010101001" => color_data <= "111111111101";
      when "000101010101010" => color_data <= "111111111101";
      when "000101010101011" => color_data <= "111111111101";
      when "000101010101100" => color_data <= "111111111101";
      when "000101010101101" => color_data <= "111111111101";
      when "000101010101110" => color_data <= "111111111101";
      when "000101010101111" => color_data <= "111111111101";
      when "000101010110000" => color_data <= "111111111101";
      when "000101010110001" => color_data <= "111111111110";
      when "000101010110010" => color_data <= "111111101000";
      when "000101010110011" => color_data <= "111111100101";
      when "000101010110100" => color_data <= "111111100111";
      when "000101010110101" => color_data <= "111111100111";
      when "000101010110110" => color_data <= "111111100111";
      when "000101010110111" => color_data <= "111111100111";
      when "000101010111000" => color_data <= "111111100111";
      when "000101010111001" => color_data <= "111111100111";
      when "000101010111010" => color_data <= "111111100111";
      when "000101010111011" => color_data <= "111111100111";
      when "000101010111100" => color_data <= "111111100111";
      when "000101010111101" => color_data <= "111111100111";
      when "000101010111110" => color_data <= "111111100111";
      when "000101010111111" => color_data <= "111111100111";
      when "000101011000000" => color_data <= "111111100111";
      when "000101011000001" => color_data <= "111111100111";
      when "000101011000010" => color_data <= "111111100111";
      when "000101011000011" => color_data <= "111111100111";
      when "000101011000100" => color_data <= "111111100110";
      when "000101011000101" => color_data <= "111111100111";
      when "000101011000110" => color_data <= "111111100111";
      when "000101011000111" => color_data <= "111111010100";
      when "000101011001000" => color_data <= "111111100101";
      when "000101011001001" => color_data <= "111111100111";
      when "000101011001010" => color_data <= "100110000010";
      when "000101011001011" => color_data <= "000100010001";
      when "000101011001100" => color_data <= "000000000000";
      when "000101011001101" => color_data <= "000000000000";
      when "000101011001110" => color_data <= "000000000000";
      when "000101011001111" => color_data <= "000000000000";
      when "000101011010000" => color_data <= "000000000000";
      when "000101011010001" => color_data <= "000000000000";
      when "000101011010010" => color_data <= "000000000000";
      when "000101011010011" => color_data <= "000000000000";
      when "000101011010100" => color_data <= "000000000000";
      when "000101011010101" => color_data <= "000000000000";
      when "000101011010110" => color_data <= "000000000000";
      when "000101011010111" => color_data <= "000000000000";
      when "000101011011000" => color_data <= "000000000000";
      when "000101011011001" => color_data <= "000000000000";
      when "000101011011010" => color_data <= "000000000000";
      when "000101011011011" => color_data <= "000000000000";
      when "000101011011100" => color_data <= "000000000000";
      when "000101011011101" => color_data <= "000000000000";
      when "000101011011110" => color_data <= "000000000000";
      when "000101011011111" => color_data <= "000000000000";
      when "000101011100000" => color_data <= "000000000000";
      when "000101011100001" => color_data <= "000000000000";
      when "000101011100010" => color_data <= "000000000000";
      when "000101011100011" => color_data <= "000000000000";
      when "000101100000000" => color_data <= "000000000000";
      when "000101100000001" => color_data <= "000000000000";
      when "000101100000010" => color_data <= "000000000000";
      when "000101100000011" => color_data <= "000000000000";
      when "000101100000100" => color_data <= "000000000000";
      when "000101100000101" => color_data <= "000000000000";
      when "000101100000110" => color_data <= "000000000000";
      when "000101100000111" => color_data <= "000000000000";
      when "000101100001000" => color_data <= "000000000000";
      when "000101100001001" => color_data <= "000000000000";
      when "000101100001010" => color_data <= "000000000000";
      when "000101100001011" => color_data <= "000000000000";
      when "000101100001100" => color_data <= "000000000000";
      when "000101100001101" => color_data <= "000000000000";
      when "000101100001110" => color_data <= "000000000000";
      when "000101100001111" => color_data <= "000000000000";
      when "000101100010000" => color_data <= "000000000000";
      when "000101100010001" => color_data <= "000000000000";
      when "000101100010010" => color_data <= "000000000000";
      when "000101100010011" => color_data <= "000000000000";
      when "000101100010100" => color_data <= "000000000000";
      when "000101100010101" => color_data <= "000000000000";
      when "000101100010110" => color_data <= "000000000000";
      when "000101100010111" => color_data <= "000000000000";
      when "000101100011000" => color_data <= "000000000000";
      when "000101100011001" => color_data <= "110110110000";
      when "000101100011010" => color_data <= "111111010000";
      when "000101100011011" => color_data <= "111111000000";
      when "000101100011100" => color_data <= "111111010000";
      when "000101100011101" => color_data <= "111111111101";
      when "000101100011110" => color_data <= "111111111110";
      when "000101100011111" => color_data <= "111111111100";
      when "000101100100000" => color_data <= "111111111101";
      when "000101100100001" => color_data <= "111111111101";
      when "000101100100010" => color_data <= "111111111101";
      when "000101100100011" => color_data <= "111111111101";
      when "000101100100100" => color_data <= "111111111101";
      when "000101100100101" => color_data <= "111111111101";
      when "000101100100110" => color_data <= "111111111101";
      when "000101100100111" => color_data <= "111111111101";
      when "000101100101000" => color_data <= "111111111101";
      when "000101100101001" => color_data <= "111111111101";
      when "000101100101010" => color_data <= "111111111101";
      when "000101100101011" => color_data <= "111111111101";
      when "000101100101100" => color_data <= "111111111101";
      when "000101100101101" => color_data <= "111111111101";
      when "000101100101110" => color_data <= "111111111101";
      when "000101100101111" => color_data <= "111111111101";
      when "000101100110000" => color_data <= "111111111101";
      when "000101100110001" => color_data <= "111111111110";
      when "000101100110010" => color_data <= "111111101000";
      when "000101100110011" => color_data <= "111111010101";
      when "000101100110100" => color_data <= "111111100111";
      when "000101100110101" => color_data <= "111111100111";
      when "000101100110110" => color_data <= "111111100111";
      when "000101100110111" => color_data <= "111111100111";
      when "000101100111000" => color_data <= "111111100111";
      when "000101100111001" => color_data <= "111111100111";
      when "000101100111010" => color_data <= "111111100111";
      when "000101100111011" => color_data <= "111111100111";
      when "000101100111100" => color_data <= "111111100111";
      when "000101100111101" => color_data <= "111111100111";
      when "000101100111110" => color_data <= "111111100111";
      when "000101100111111" => color_data <= "111111100111";
      when "000101101000000" => color_data <= "111111100111";
      when "000101101000001" => color_data <= "111111100111";
      when "000101101000010" => color_data <= "111111100111";
      when "000101101000011" => color_data <= "111111100111";
      when "000101101000100" => color_data <= "111111100111";
      when "000101101000101" => color_data <= "111111100110";
      when "000101101000110" => color_data <= "111111100111";
      when "000101101000111" => color_data <= "111111100111";
      when "000101101001000" => color_data <= "111111010100";
      when "000101101001001" => color_data <= "111111100110";
      when "000101101001010" => color_data <= "111111010100";
      when "000101101001011" => color_data <= "100110000010";
      when "000101101001100" => color_data <= "000000000000";
      when "000101101001101" => color_data <= "000000000000";
      when "000101101001110" => color_data <= "000000000000";
      when "000101101001111" => color_data <= "000000000000";
      when "000101101010000" => color_data <= "000000000000";
      when "000101101010001" => color_data <= "000000000000";
      when "000101101010010" => color_data <= "000000000000";
      when "000101101010011" => color_data <= "000000000000";
      when "000101101010100" => color_data <= "000000000000";
      when "000101101010101" => color_data <= "000000000000";
      when "000101101010110" => color_data <= "000000000000";
      when "000101101010111" => color_data <= "000000000000";
      when "000101101011000" => color_data <= "000000000000";
      when "000101101011001" => color_data <= "000000000000";
      when "000101101011010" => color_data <= "000000000000";
      when "000101101011011" => color_data <= "000000000000";
      when "000101101011100" => color_data <= "000000000000";
      when "000101101011101" => color_data <= "000000000000";
      when "000101101011110" => color_data <= "000000000000";
      when "000101101011111" => color_data <= "000000000000";
      when "000101101100000" => color_data <= "000000000000";
      when "000101101100001" => color_data <= "000000000000";
      when "000101101100010" => color_data <= "000000000000";
      when "000101101100011" => color_data <= "000000000000";
      when "000101110000000" => color_data <= "000000000000";
      when "000101110000001" => color_data <= "000000000000";
      when "000101110000010" => color_data <= "000000000000";
      when "000101110000011" => color_data <= "000000000000";
      when "000101110000100" => color_data <= "000000000000";
      when "000101110000101" => color_data <= "000000000000";
      when "000101110000110" => color_data <= "000000000000";
      when "000101110000111" => color_data <= "000000000000";
      when "000101110001000" => color_data <= "000000000000";
      when "000101110001001" => color_data <= "000000000000";
      when "000101110001010" => color_data <= "000000000000";
      when "000101110001011" => color_data <= "000000000000";
      when "000101110001100" => color_data <= "000000000000";
      when "000101110001101" => color_data <= "000000000000";
      when "000101110001110" => color_data <= "000000000000";
      when "000101110001111" => color_data <= "000000000000";
      when "000101110010000" => color_data <= "000000000000";
      when "000101110010001" => color_data <= "000000000000";
      when "000101110010010" => color_data <= "000000000000";
      when "000101110010011" => color_data <= "000000000000";
      when "000101110010100" => color_data <= "000000000000";
      when "000101110010101" => color_data <= "000000000000";
      when "000101110010110" => color_data <= "000000000000";
      when "000101110010111" => color_data <= "000000000000";
      when "000101110011000" => color_data <= "101010010010";
      when "000101110011001" => color_data <= "111111000000";
      when "000101110011010" => color_data <= "111111010001";
      when "000101110011011" => color_data <= "111111000000";
      when "000101110011100" => color_data <= "111111100110";
      when "000101110011101" => color_data <= "111111111111";
      when "000101110011110" => color_data <= "111111111100";
      when "000101110011111" => color_data <= "111111111101";
      when "000101110100000" => color_data <= "111111111101";
      when "000101110100001" => color_data <= "111111111101";
      when "000101110100010" => color_data <= "111111111101";
      when "000101110100011" => color_data <= "111111111101";
      when "000101110100100" => color_data <= "111111111101";
      when "000101110100101" => color_data <= "111111111101";
      when "000101110100110" => color_data <= "111111111101";
      when "000101110100111" => color_data <= "111111111101";
      when "000101110101000" => color_data <= "111111111101";
      when "000101110101001" => color_data <= "111111111101";
      when "000101110101010" => color_data <= "111111111101";
      when "000101110101011" => color_data <= "111111111101";
      when "000101110101100" => color_data <= "111111111101";
      when "000101110101101" => color_data <= "111111111101";
      when "000101110101110" => color_data <= "111111111101";
      when "000101110101111" => color_data <= "111111111101";
      when "000101110110000" => color_data <= "111111111101";
      when "000101110110001" => color_data <= "111111111110";
      when "000101110110010" => color_data <= "111111101000";
      when "000101110110011" => color_data <= "111111100101";
      when "000101110110100" => color_data <= "111111100111";
      when "000101110110101" => color_data <= "111111100111";
      when "000101110110110" => color_data <= "111111100111";
      when "000101110110111" => color_data <= "111111100111";
      when "000101110111000" => color_data <= "111111100111";
      when "000101110111001" => color_data <= "111111100111";
      when "000101110111010" => color_data <= "111111100111";
      when "000101110111011" => color_data <= "111111100111";
      when "000101110111100" => color_data <= "111111100111";
      when "000101110111101" => color_data <= "111111100111";
      when "000101110111110" => color_data <= "111111100111";
      when "000101110111111" => color_data <= "111111100111";
      when "000101111000000" => color_data <= "111111100111";
      when "000101111000001" => color_data <= "111111100111";
      when "000101111000010" => color_data <= "111111100111";
      when "000101111000011" => color_data <= "111111100111";
      when "000101111000100" => color_data <= "111111100111";
      when "000101111000101" => color_data <= "111111100111";
      when "000101111000110" => color_data <= "111111100110";
      when "000101111000111" => color_data <= "111111100111";
      when "000101111001000" => color_data <= "111111100111";
      when "000101111001001" => color_data <= "111111010010";
      when "000101111001010" => color_data <= "111111010000";
      when "000101111001011" => color_data <= "110110110000";
      when "000101111001100" => color_data <= "010101010011";
      when "000101111001101" => color_data <= "000000000000";
      when "000101111001110" => color_data <= "000000000000";
      when "000101111001111" => color_data <= "000000000000";
      when "000101111010000" => color_data <= "000000000000";
      when "000101111010001" => color_data <= "000000000000";
      when "000101111010010" => color_data <= "000000000000";
      when "000101111010011" => color_data <= "000000000000";
      when "000101111010100" => color_data <= "000000000000";
      when "000101111010101" => color_data <= "000000000000";
      when "000101111010110" => color_data <= "000000000000";
      when "000101111010111" => color_data <= "000000000000";
      when "000101111011000" => color_data <= "000000000000";
      when "000101111011001" => color_data <= "000000000000";
      when "000101111011010" => color_data <= "000000000000";
      when "000101111011011" => color_data <= "000000000000";
      when "000101111011100" => color_data <= "000000000000";
      when "000101111011101" => color_data <= "000000000000";
      when "000101111011110" => color_data <= "000000000000";
      when "000101111011111" => color_data <= "000000000000";
      when "000101111100000" => color_data <= "000000000000";
      when "000101111100001" => color_data <= "000000000000";
      when "000101111100010" => color_data <= "000000000000";
      when "000101111100011" => color_data <= "000000000000";
      when "000110000000000" => color_data <= "000000000000";
      when "000110000000001" => color_data <= "000000000000";
      when "000110000000010" => color_data <= "000000000000";
      when "000110000000011" => color_data <= "000000000000";
      when "000110000000100" => color_data <= "000000000000";
      when "000110000000101" => color_data <= "000000000000";
      when "000110000000110" => color_data <= "000000000000";
      when "000110000000111" => color_data <= "000000000000";
      when "000110000001000" => color_data <= "000000000000";
      when "000110000001001" => color_data <= "000000000000";
      when "000110000001010" => color_data <= "000000000000";
      when "000110000001011" => color_data <= "000000000000";
      when "000110000001100" => color_data <= "000000000000";
      when "000110000001101" => color_data <= "000000000000";
      when "000110000001110" => color_data <= "000000000000";
      when "000110000001111" => color_data <= "000000000000";
      when "000110000010000" => color_data <= "000000000000";
      when "000110000010001" => color_data <= "000000000000";
      when "000110000010010" => color_data <= "000000000000";
      when "000110000010011" => color_data <= "000000000000";
      when "000110000010100" => color_data <= "000000000000";
      when "000110000010101" => color_data <= "000000000000";
      when "000110000010110" => color_data <= "000000000000";
      when "000110000010111" => color_data <= "001000100001";
      when "000110000011000" => color_data <= "110110110000";
      when "000110000011001" => color_data <= "111111010000";
      when "000110000011010" => color_data <= "111111010000";
      when "000110000011011" => color_data <= "111111000000";
      when "000110000011100" => color_data <= "111111101001";
      when "000110000011101" => color_data <= "111111111111";
      when "000110000011110" => color_data <= "111111111101";
      when "000110000011111" => color_data <= "111111111101";
      when "000110000100000" => color_data <= "111111111100";
      when "000110000100001" => color_data <= "111111111101";
      when "000110000100010" => color_data <= "111111111101";
      when "000110000100011" => color_data <= "111111111101";
      when "000110000100100" => color_data <= "111111111101";
      when "000110000100101" => color_data <= "111111111101";
      when "000110000100110" => color_data <= "111111111101";
      when "000110000100111" => color_data <= "111111111101";
      when "000110000101000" => color_data <= "111111111101";
      when "000110000101001" => color_data <= "111111111101";
      when "000110000101010" => color_data <= "111111111101";
      when "000110000101011" => color_data <= "111111111101";
      when "000110000101100" => color_data <= "111111111101";
      when "000110000101101" => color_data <= "111111111101";
      when "000110000101110" => color_data <= "111111111101";
      when "000110000101111" => color_data <= "111111111101";
      when "000110000110000" => color_data <= "111111111101";
      when "000110000110001" => color_data <= "111111111110";
      when "000110000110010" => color_data <= "111111100111";
      when "000110000110011" => color_data <= "111111100101";
      when "000110000110100" => color_data <= "111111100111";
      when "000110000110101" => color_data <= "111111100111";
      when "000110000110110" => color_data <= "111111100111";
      when "000110000110111" => color_data <= "111111100111";
      when "000110000111000" => color_data <= "111111100111";
      when "000110000111001" => color_data <= "111111100111";
      when "000110000111010" => color_data <= "111111100111";
      when "000110000111011" => color_data <= "111111100111";
      when "000110000111100" => color_data <= "111111100111";
      when "000110000111101" => color_data <= "111111100111";
      when "000110000111110" => color_data <= "111111100111";
      when "000110000111111" => color_data <= "111111100111";
      when "000110001000000" => color_data <= "111111100111";
      when "000110001000001" => color_data <= "111111100111";
      when "000110001000010" => color_data <= "111111100111";
      when "000110001000011" => color_data <= "111111100111";
      when "000110001000100" => color_data <= "111111100111";
      when "000110001000101" => color_data <= "111111100110";
      when "000110001000110" => color_data <= "111111100110";
      when "000110001000111" => color_data <= "111111100111";
      when "000110001001000" => color_data <= "111111101000";
      when "000110001001001" => color_data <= "111111010100";
      when "000110001001010" => color_data <= "111111010000";
      when "000110001001011" => color_data <= "111111010000";
      when "000110001001100" => color_data <= "110110110000";
      when "000110001001101" => color_data <= "000000000000";
      when "000110001001110" => color_data <= "000000000000";
      when "000110001001111" => color_data <= "000000000000";
      when "000110001010000" => color_data <= "000000000000";
      when "000110001010001" => color_data <= "000000000000";
      when "000110001010010" => color_data <= "000000000000";
      when "000110001010011" => color_data <= "000000000000";
      when "000110001010100" => color_data <= "000000000000";
      when "000110001010101" => color_data <= "000000000000";
      when "000110001010110" => color_data <= "000000000000";
      when "000110001010111" => color_data <= "000000000000";
      when "000110001011000" => color_data <= "000000000000";
      when "000110001011001" => color_data <= "000000000000";
      when "000110001011010" => color_data <= "000000000000";
      when "000110001011011" => color_data <= "000000000000";
      when "000110001011100" => color_data <= "000000000000";
      when "000110001011101" => color_data <= "000000000000";
      when "000110001011110" => color_data <= "000000000000";
      when "000110001011111" => color_data <= "000000000000";
      when "000110001100000" => color_data <= "000000000000";
      when "000110001100001" => color_data <= "000000000000";
      when "000110001100010" => color_data <= "000000000000";
      when "000110001100011" => color_data <= "000000000000";
      when "000110010000000" => color_data <= "000000000000";
      when "000110010000001" => color_data <= "000000000000";
      when "000110010000010" => color_data <= "000000000000";
      when "000110010000011" => color_data <= "000000000000";
      when "000110010000100" => color_data <= "000000000000";
      when "000110010000101" => color_data <= "000000000000";
      when "000110010000110" => color_data <= "000000000000";
      when "000110010000111" => color_data <= "000000000000";
      when "000110010001000" => color_data <= "000000000000";
      when "000110010001001" => color_data <= "000000000000";
      when "000110010001010" => color_data <= "000000000000";
      when "000110010001011" => color_data <= "000000000000";
      when "000110010001100" => color_data <= "000000000000";
      when "000110010001101" => color_data <= "000000000000";
      when "000110010001110" => color_data <= "000000000000";
      when "000110010001111" => color_data <= "000000000000";
      when "000110010010000" => color_data <= "000000000000";
      when "000110010010001" => color_data <= "000000000000";
      when "000110010010010" => color_data <= "000000000000";
      when "000110010010011" => color_data <= "000000000000";
      when "000110010010100" => color_data <= "000000000000";
      when "000110010010101" => color_data <= "000000000000";
      when "000110010010110" => color_data <= "000000000000";
      when "000110010010111" => color_data <= "101010010010";
      when "000110010011000" => color_data <= "111111000000";
      when "000110010011001" => color_data <= "111111010001";
      when "000110010011010" => color_data <= "111111010000";
      when "000110010011011" => color_data <= "111111010000";
      when "000110010011100" => color_data <= "111111111011";
      when "000110010011101" => color_data <= "111111111110";
      when "000110010011110" => color_data <= "111111111101";
      when "000110010011111" => color_data <= "111111111101";
      when "000110010100000" => color_data <= "111111111101";
      when "000110010100001" => color_data <= "111111111101";
      when "000110010100010" => color_data <= "111111111101";
      when "000110010100011" => color_data <= "111111111101";
      when "000110010100100" => color_data <= "111111111101";
      when "000110010100101" => color_data <= "111111111101";
      when "000110010100110" => color_data <= "111111111101";
      when "000110010100111" => color_data <= "111111111101";
      when "000110010101000" => color_data <= "111111111101";
      when "000110010101001" => color_data <= "111111111101";
      when "000110010101010" => color_data <= "111111111101";
      when "000110010101011" => color_data <= "111111111101";
      when "000110010101100" => color_data <= "111111111101";
      when "000110010101101" => color_data <= "111111111101";
      when "000110010101110" => color_data <= "111111111101";
      when "000110010101111" => color_data <= "111111111101";
      when "000110010110000" => color_data <= "111111111101";
      when "000110010110001" => color_data <= "111111111110";
      when "000110010110010" => color_data <= "111111100111";
      when "000110010110011" => color_data <= "111111100101";
      when "000110010110100" => color_data <= "111111100111";
      when "000110010110101" => color_data <= "111111100111";
      when "000110010110110" => color_data <= "111111100111";
      when "000110010110111" => color_data <= "111111100111";
      when "000110010111000" => color_data <= "111111100111";
      when "000110010111001" => color_data <= "111111100111";
      when "000110010111010" => color_data <= "111111100111";
      when "000110010111011" => color_data <= "111111100111";
      when "000110010111100" => color_data <= "111111100111";
      when "000110010111101" => color_data <= "111111100111";
      when "000110010111110" => color_data <= "111111100111";
      when "000110010111111" => color_data <= "111111100111";
      when "000110011000000" => color_data <= "111111100111";
      when "000110011000001" => color_data <= "111111100111";
      when "000110011000010" => color_data <= "111111100111";
      when "000110011000011" => color_data <= "111111100111";
      when "000110011000100" => color_data <= "111111100110";
      when "000110011000101" => color_data <= "111111100111";
      when "000110011000110" => color_data <= "111111100111";
      when "000110011000111" => color_data <= "111111100110";
      when "000110011001000" => color_data <= "111111100111";
      when "000110011001001" => color_data <= "111111100101";
      when "000110011001010" => color_data <= "111111010000";
      when "000110011001011" => color_data <= "111111010000";
      when "000110011001100" => color_data <= "111111000000";
      when "000110011001101" => color_data <= "011101100011";
      when "000110011001110" => color_data <= "000000000000";
      when "000110011001111" => color_data <= "000000000000";
      when "000110011010000" => color_data <= "000000000000";
      when "000110011010001" => color_data <= "000000000000";
      when "000110011010010" => color_data <= "000000000000";
      when "000110011010011" => color_data <= "000000000000";
      when "000110011010100" => color_data <= "000000000000";
      when "000110011010101" => color_data <= "000000000000";
      when "000110011010110" => color_data <= "000000000000";
      when "000110011010111" => color_data <= "000000000000";
      when "000110011011000" => color_data <= "000000000000";
      when "000110011011001" => color_data <= "000000000000";
      when "000110011011010" => color_data <= "000000000000";
      when "000110011011011" => color_data <= "000000000000";
      when "000110011011100" => color_data <= "000000000000";
      when "000110011011101" => color_data <= "000000000000";
      when "000110011011110" => color_data <= "000000000000";
      when "000110011011111" => color_data <= "000000000000";
      when "000110011100000" => color_data <= "000000000000";
      when "000110011100001" => color_data <= "000000000000";
      when "000110011100010" => color_data <= "000000000000";
      when "000110011100011" => color_data <= "000000000000";
      when "000110100000000" => color_data <= "000000000000";
      when "000110100000001" => color_data <= "000000000000";
      when "000110100000010" => color_data <= "000000000000";
      when "000110100000011" => color_data <= "000000000000";
      when "000110100000100" => color_data <= "000000000000";
      when "000110100000101" => color_data <= "000000000000";
      when "000110100000110" => color_data <= "000000000000";
      when "000110100000111" => color_data <= "000000000000";
      when "000110100001000" => color_data <= "000000000000";
      when "000110100001001" => color_data <= "000000000000";
      when "000110100001010" => color_data <= "000000000000";
      when "000110100001011" => color_data <= "000000000000";
      when "000110100001100" => color_data <= "000000000000";
      when "000110100001101" => color_data <= "000000000000";
      when "000110100001110" => color_data <= "000000000000";
      when "000110100001111" => color_data <= "000000000000";
      when "000110100010000" => color_data <= "000000000000";
      when "000110100010001" => color_data <= "000000000000";
      when "000110100010010" => color_data <= "000000000000";
      when "000110100010011" => color_data <= "000000000000";
      when "000110100010100" => color_data <= "000000000000";
      when "000110100010101" => color_data <= "000000000000";
      when "000110100010110" => color_data <= "001000100001";
      when "000110100010111" => color_data <= "110110110000";
      when "000110100011000" => color_data <= "111111010000";
      when "000110100011001" => color_data <= "111111010000";
      when "000110100011010" => color_data <= "111111010000";
      when "000110100011011" => color_data <= "111111010010";
      when "000110100011100" => color_data <= "111111111100";
      when "000110100011101" => color_data <= "111111111101";
      when "000110100011110" => color_data <= "111111111100";
      when "000110100011111" => color_data <= "111111111101";
      when "000110100100000" => color_data <= "111111111110";
      when "000110100100001" => color_data <= "111111111101";
      when "000110100100010" => color_data <= "111111111100";
      when "000110100100011" => color_data <= "111111111101";
      when "000110100100100" => color_data <= "111111111101";
      when "000110100100101" => color_data <= "111111111101";
      when "000110100100110" => color_data <= "111111111101";
      when "000110100100111" => color_data <= "111111111101";
      when "000110100101000" => color_data <= "111111111101";
      when "000110100101001" => color_data <= "111111111101";
      when "000110100101010" => color_data <= "111111111101";
      when "000110100101011" => color_data <= "111111111101";
      when "000110100101100" => color_data <= "111111111101";
      when "000110100101101" => color_data <= "111111111101";
      when "000110100101110" => color_data <= "111111111101";
      when "000110100101111" => color_data <= "111111111101";
      when "000110100110000" => color_data <= "111111111101";
      when "000110100110001" => color_data <= "111111111110";
      when "000110100110010" => color_data <= "111111100111";
      when "000110100110011" => color_data <= "111111100101";
      when "000110100110100" => color_data <= "111111100111";
      when "000110100110101" => color_data <= "111111100111";
      when "000110100110110" => color_data <= "111111100111";
      when "000110100110111" => color_data <= "111111100111";
      when "000110100111000" => color_data <= "111111100111";
      when "000110100111001" => color_data <= "111111100111";
      when "000110100111010" => color_data <= "111111100111";
      when "000110100111011" => color_data <= "111111100111";
      when "000110100111100" => color_data <= "111111100111";
      when "000110100111101" => color_data <= "111111100111";
      when "000110100111110" => color_data <= "111111100111";
      when "000110100111111" => color_data <= "111111100111";
      when "000110101000000" => color_data <= "111111100111";
      when "000110101000001" => color_data <= "111111100111";
      when "000110101000010" => color_data <= "111111100111";
      when "000110101000011" => color_data <= "111111100111";
      when "000110101000100" => color_data <= "111111100110";
      when "000110101000101" => color_data <= "111111101000";
      when "000110101000110" => color_data <= "111111111011";
      when "000110101000111" => color_data <= "111111101000";
      when "000110101001000" => color_data <= "111111100110";
      when "000110101001001" => color_data <= "111111100110";
      when "000110101001010" => color_data <= "111111010001";
      when "000110101001011" => color_data <= "111111010000";
      when "000110101001100" => color_data <= "111111010000";
      when "000110101001101" => color_data <= "110010110000";
      when "000110101001110" => color_data <= "000000000000";
      when "000110101001111" => color_data <= "000000000000";
      when "000110101010000" => color_data <= "000000000000";
      when "000110101010001" => color_data <= "000000000000";
      when "000110101010010" => color_data <= "000000000000";
      when "000110101010011" => color_data <= "000000000000";
      when "000110101010100" => color_data <= "000000000000";
      when "000110101010101" => color_data <= "000000000000";
      when "000110101010110" => color_data <= "000000000000";
      when "000110101010111" => color_data <= "000000000000";
      when "000110101011000" => color_data <= "000000000000";
      when "000110101011001" => color_data <= "000000000000";
      when "000110101011010" => color_data <= "000000000000";
      when "000110101011011" => color_data <= "000000000000";
      when "000110101011100" => color_data <= "000000000000";
      when "000110101011101" => color_data <= "000000000000";
      when "000110101011110" => color_data <= "000000000000";
      when "000110101011111" => color_data <= "000000000000";
      when "000110101100000" => color_data <= "000000000000";
      when "000110101100001" => color_data <= "000000000000";
      when "000110101100010" => color_data <= "000000000000";
      when "000110101100011" => color_data <= "000000000000";
      when "000110110000000" => color_data <= "000000000000";
      when "000110110000001" => color_data <= "000000000000";
      when "000110110000010" => color_data <= "000000000000";
      when "000110110000011" => color_data <= "000000000000";
      when "000110110000100" => color_data <= "000000000000";
      when "000110110000101" => color_data <= "000000000000";
      when "000110110000110" => color_data <= "000000000000";
      when "000110110000111" => color_data <= "000000000000";
      when "000110110001000" => color_data <= "000000000000";
      when "000110110001001" => color_data <= "000000000000";
      when "000110110001010" => color_data <= "000000000000";
      when "000110110001011" => color_data <= "000000000000";
      when "000110110001100" => color_data <= "000000000000";
      when "000110110001101" => color_data <= "000000000000";
      when "000110110001110" => color_data <= "000000000000";
      when "000110110001111" => color_data <= "000000000000";
      when "000110110010000" => color_data <= "000000000000";
      when "000110110010001" => color_data <= "000000000000";
      when "000110110010010" => color_data <= "000000000000";
      when "000110110010011" => color_data <= "000000000000";
      when "000110110010100" => color_data <= "000000000000";
      when "000110110010101" => color_data <= "000000000000";
      when "000110110010110" => color_data <= "100110000010";
      when "000110110010111" => color_data <= "111111000000";
      when "000110110011000" => color_data <= "111111010000";
      when "000110110011001" => color_data <= "111111010000";
      when "000110110011010" => color_data <= "111111000000";
      when "000110110011011" => color_data <= "111111010010";
      when "000110110011100" => color_data <= "111111111101";
      when "000110110011101" => color_data <= "111111111101";
      when "000110110011110" => color_data <= "111111111100";
      when "000110110011111" => color_data <= "111111111101";
      when "000110110100000" => color_data <= "111111111110";
      when "000110110100001" => color_data <= "111111111101";
      when "000110110100010" => color_data <= "111111111100";
      when "000110110100011" => color_data <= "111111111101";
      when "000110110100100" => color_data <= "111111111101";
      when "000110110100101" => color_data <= "111111111101";
      when "000110110100110" => color_data <= "111111111101";
      when "000110110100111" => color_data <= "111111111101";
      when "000110110101000" => color_data <= "111111111101";
      when "000110110101001" => color_data <= "111111111101";
      when "000110110101010" => color_data <= "111111111101";
      when "000110110101011" => color_data <= "111111111101";
      when "000110110101100" => color_data <= "111111111101";
      when "000110110101101" => color_data <= "111111111101";
      when "000110110101110" => color_data <= "111111111101";
      when "000110110101111" => color_data <= "111111111101";
      when "000110110110000" => color_data <= "111111111101";
      when "000110110110001" => color_data <= "111111111110";
      when "000110110110010" => color_data <= "111111100111";
      when "000110110110011" => color_data <= "111111100101";
      when "000110110110100" => color_data <= "111111100111";
      when "000110110110101" => color_data <= "111111100111";
      when "000110110110110" => color_data <= "111111100111";
      when "000110110110111" => color_data <= "111111100111";
      when "000110110111000" => color_data <= "111111100111";
      when "000110110111001" => color_data <= "111111100111";
      when "000110110111010" => color_data <= "111111100111";
      when "000110110111011" => color_data <= "111111100111";
      when "000110110111100" => color_data <= "111111100111";
      when "000110110111101" => color_data <= "111111100111";
      when "000110110111110" => color_data <= "111111100111";
      when "000110110111111" => color_data <= "111111100111";
      when "000110111000000" => color_data <= "111111100111";
      when "000110111000001" => color_data <= "111111100111";
      when "000110111000010" => color_data <= "111111100111";
      when "000110111000011" => color_data <= "111111100111";
      when "000110111000100" => color_data <= "111111100110";
      when "000110111000101" => color_data <= "111111101000";
      when "000110111000110" => color_data <= "111111111011";
      when "000110111000111" => color_data <= "111111101000";
      when "000110111001000" => color_data <= "111111100110";
      when "000110111001001" => color_data <= "111111100111";
      when "000110111001010" => color_data <= "111111010010";
      when "000110111001011" => color_data <= "111111010000";
      when "000110111001100" => color_data <= "111111010000";
      when "000110111001101" => color_data <= "110110110000";
      when "000110111001110" => color_data <= "010101010011";
      when "000110111001111" => color_data <= "000000000000";
      when "000110111010000" => color_data <= "000000000000";
      when "000110111010001" => color_data <= "000000000000";
      when "000110111010010" => color_data <= "000000000000";
      when "000110111010011" => color_data <= "000000000000";
      when "000110111010100" => color_data <= "000000000000";
      when "000110111010101" => color_data <= "000000000000";
      when "000110111010110" => color_data <= "000000000000";
      when "000110111010111" => color_data <= "000000000000";
      when "000110111011000" => color_data <= "000000000000";
      when "000110111011001" => color_data <= "000000000000";
      when "000110111011010" => color_data <= "000000000000";
      when "000110111011011" => color_data <= "000000000000";
      when "000110111011100" => color_data <= "000000000000";
      when "000110111011101" => color_data <= "000000000000";
      when "000110111011110" => color_data <= "000000000000";
      when "000110111011111" => color_data <= "000000000000";
      when "000110111100000" => color_data <= "000000000000";
      when "000110111100001" => color_data <= "000000000000";
      when "000110111100010" => color_data <= "000000000000";
      when "000110111100011" => color_data <= "000000000000";
      when "000111000000000" => color_data <= "000000000000";
      when "000111000000001" => color_data <= "000000000000";
      when "000111000000010" => color_data <= "000000000000";
      when "000111000000011" => color_data <= "000000000000";
      when "000111000000100" => color_data <= "000000000000";
      when "000111000000101" => color_data <= "000000000000";
      when "000111000000110" => color_data <= "000000000000";
      when "000111000000111" => color_data <= "000000000000";
      when "000111000001000" => color_data <= "000000000000";
      when "000111000001001" => color_data <= "000000000000";
      when "000111000001010" => color_data <= "000000000000";
      when "000111000001011" => color_data <= "000000000000";
      when "000111000001100" => color_data <= "000000000000";
      when "000111000001101" => color_data <= "000000000000";
      when "000111000001110" => color_data <= "000000000000";
      when "000111000001111" => color_data <= "000000000000";
      when "000111000010000" => color_data <= "000000000000";
      when "000111000010001" => color_data <= "000000000000";
      when "000111000010010" => color_data <= "000000000000";
      when "000111000010011" => color_data <= "000000000000";
      when "000111000010100" => color_data <= "000000000000";
      when "000111000010101" => color_data <= "000000000000";
      when "000111000010110" => color_data <= "110110110000";
      when "000111000010111" => color_data <= "111111010000";
      when "000111000011000" => color_data <= "111111010000";
      when "000111000011001" => color_data <= "111111010000";
      when "000111000011010" => color_data <= "111111010000";
      when "000111000011011" => color_data <= "111111010010";
      when "000111000011100" => color_data <= "111111111101";
      when "000111000011101" => color_data <= "111111111101";
      when "000111000011110" => color_data <= "111111111100";
      when "000111000011111" => color_data <= "111111111101";
      when "000111000100000" => color_data <= "111111111110";
      when "000111000100001" => color_data <= "111111111101";
      when "000111000100010" => color_data <= "111111111100";
      when "000111000100011" => color_data <= "111111111101";
      when "000111000100100" => color_data <= "111111111101";
      when "000111000100101" => color_data <= "111111111101";
      when "000111000100110" => color_data <= "111111111101";
      when "000111000100111" => color_data <= "111111111101";
      when "000111000101000" => color_data <= "111111111101";
      when "000111000101001" => color_data <= "111111111101";
      when "000111000101010" => color_data <= "111111111101";
      when "000111000101011" => color_data <= "111111111101";
      when "000111000101100" => color_data <= "111111111101";
      when "000111000101101" => color_data <= "111111111101";
      when "000111000101110" => color_data <= "111111111101";
      when "000111000101111" => color_data <= "111111111101";
      when "000111000110000" => color_data <= "111111111101";
      when "000111000110001" => color_data <= "111111111110";
      when "000111000110010" => color_data <= "111111101000";
      when "000111000110011" => color_data <= "111111100101";
      when "000111000110100" => color_data <= "111111100111";
      when "000111000110101" => color_data <= "111111100111";
      when "000111000110110" => color_data <= "111111100111";
      when "000111000110111" => color_data <= "111111100111";
      when "000111000111000" => color_data <= "111111100111";
      when "000111000111001" => color_data <= "111111100111";
      when "000111000111010" => color_data <= "111111100111";
      when "000111000111011" => color_data <= "111111100111";
      when "000111000111100" => color_data <= "111111100111";
      when "000111000111101" => color_data <= "111111100111";
      when "000111000111110" => color_data <= "111111100111";
      when "000111000111111" => color_data <= "111111100111";
      when "000111001000000" => color_data <= "111111100111";
      when "000111001000001" => color_data <= "111111100111";
      when "000111001000010" => color_data <= "111111100111";
      when "000111001000011" => color_data <= "111111100111";
      when "000111001000100" => color_data <= "111111100110";
      when "000111001000101" => color_data <= "111111101000";
      when "000111001000110" => color_data <= "111111111011";
      when "000111001000111" => color_data <= "111111101000";
      when "000111001001000" => color_data <= "111111100110";
      when "000111001001001" => color_data <= "111111100111";
      when "000111001001010" => color_data <= "111111010010";
      when "000111001001011" => color_data <= "111111010000";
      when "000111001001100" => color_data <= "111111010001";
      when "000111001001101" => color_data <= "111111010000";
      when "000111001001110" => color_data <= "101110010001";
      when "000111001001111" => color_data <= "000000000000";
      when "000111001010000" => color_data <= "000000000000";
      when "000111001010001" => color_data <= "000000000000";
      when "000111001010010" => color_data <= "000000000000";
      when "000111001010011" => color_data <= "000000000000";
      when "000111001010100" => color_data <= "000000000000";
      when "000111001010101" => color_data <= "000000000000";
      when "000111001010110" => color_data <= "000000000000";
      when "000111001010111" => color_data <= "000000000000";
      when "000111001011000" => color_data <= "000000000000";
      when "000111001011001" => color_data <= "000000000000";
      when "000111001011010" => color_data <= "000000000000";
      when "000111001011011" => color_data <= "000000000000";
      when "000111001011100" => color_data <= "000000000000";
      when "000111001011101" => color_data <= "000000000000";
      when "000111001011110" => color_data <= "000000000000";
      when "000111001011111" => color_data <= "000000000000";
      when "000111001100000" => color_data <= "000000000000";
      when "000111001100001" => color_data <= "000000000000";
      when "000111001100010" => color_data <= "000000000000";
      when "000111001100011" => color_data <= "000000000000";
      when "000111010000000" => color_data <= "000000000000";
      when "000111010000001" => color_data <= "000000000000";
      when "000111010000010" => color_data <= "000000000000";
      when "000111010000011" => color_data <= "000000000000";
      when "000111010000100" => color_data <= "000000000000";
      when "000111010000101" => color_data <= "000000000000";
      when "000111010000110" => color_data <= "000000000000";
      when "000111010000111" => color_data <= "000000000000";
      when "000111010001000" => color_data <= "000000000000";
      when "000111010001001" => color_data <= "000000000000";
      when "000111010001010" => color_data <= "000000000000";
      when "000111010001011" => color_data <= "000000000000";
      when "000111010001100" => color_data <= "000000000000";
      when "000111010001101" => color_data <= "000000000000";
      when "000111010001110" => color_data <= "000000000000";
      when "000111010001111" => color_data <= "000000000000";
      when "000111010010000" => color_data <= "000000000000";
      when "000111010010001" => color_data <= "000000000000";
      when "000111010010010" => color_data <= "000000000000";
      when "000111010010011" => color_data <= "000000000000";
      when "000111010010100" => color_data <= "000000000000";
      when "000111010010101" => color_data <= "010101010011";
      when "000111010010110" => color_data <= "111111000000";
      when "000111010010111" => color_data <= "111111010000";
      when "000111010011000" => color_data <= "111111010000";
      when "000111010011001" => color_data <= "111111010000";
      when "000111010011010" => color_data <= "111111010000";
      when "000111010011011" => color_data <= "111111010011";
      when "000111010011100" => color_data <= "111111111101";
      when "000111010011101" => color_data <= "111111111101";
      when "000111010011110" => color_data <= "111111111101";
      when "000111010011111" => color_data <= "111111111101";
      when "000111010100000" => color_data <= "111111111101";
      when "000111010100001" => color_data <= "111111111100";
      when "000111010100010" => color_data <= "111111111100";
      when "000111010100011" => color_data <= "111111111101";
      when "000111010100100" => color_data <= "111111111101";
      when "000111010100101" => color_data <= "111111111101";
      when "000111010100110" => color_data <= "111111111101";
      when "000111010100111" => color_data <= "111111111101";
      when "000111010101000" => color_data <= "111111111101";
      when "000111010101001" => color_data <= "111111111101";
      when "000111010101010" => color_data <= "111111111101";
      when "000111010101011" => color_data <= "111111111101";
      when "000111010101100" => color_data <= "111111111101";
      when "000111010101101" => color_data <= "111111111101";
      when "000111010101110" => color_data <= "111111111101";
      when "000111010101111" => color_data <= "111111111101";
      when "000111010110000" => color_data <= "111111111101";
      when "000111010110001" => color_data <= "111111111101";
      when "000111010110010" => color_data <= "111111101000";
      when "000111010110011" => color_data <= "111111100101";
      when "000111010110100" => color_data <= "111111100111";
      when "000111010110101" => color_data <= "111111100111";
      when "000111010110110" => color_data <= "111111100111";
      when "000111010110111" => color_data <= "111111100111";
      when "000111010111000" => color_data <= "111111100111";
      when "000111010111001" => color_data <= "111111100111";
      when "000111010111010" => color_data <= "111111100111";
      when "000111010111011" => color_data <= "111111100111";
      when "000111010111100" => color_data <= "111111100111";
      when "000111010111101" => color_data <= "111111100111";
      when "000111010111110" => color_data <= "111111100111";
      when "000111010111111" => color_data <= "111111100111";
      when "000111011000000" => color_data <= "111111100111";
      when "000111011000001" => color_data <= "111111100111";
      when "000111011000010" => color_data <= "111111100111";
      when "000111011000011" => color_data <= "111111100111";
      when "000111011000100" => color_data <= "111111100110";
      when "000111011000101" => color_data <= "111111100111";
      when "000111011000110" => color_data <= "111111100111";
      when "000111011000111" => color_data <= "111111100111";
      when "000111011001000" => color_data <= "111111100111";
      when "000111011001001" => color_data <= "111111100111";
      when "000111011001010" => color_data <= "111111010011";
      when "000111011001011" => color_data <= "111111010000";
      when "000111011001100" => color_data <= "111111010000";
      when "000111011001101" => color_data <= "111111010000";
      when "000111011001110" => color_data <= "110110110000";
      when "000111011001111" => color_data <= "001000100001";
      when "000111011010000" => color_data <= "000000000000";
      when "000111011010001" => color_data <= "000000000000";
      when "000111011010010" => color_data <= "000000000000";
      when "000111011010011" => color_data <= "000000000000";
      when "000111011010100" => color_data <= "000000000000";
      when "000111011010101" => color_data <= "000000000000";
      when "000111011010110" => color_data <= "000000000000";
      when "000111011010111" => color_data <= "000000000000";
      when "000111011011000" => color_data <= "000000000000";
      when "000111011011001" => color_data <= "000000000000";
      when "000111011011010" => color_data <= "000000000000";
      when "000111011011011" => color_data <= "000000000000";
      when "000111011011100" => color_data <= "000000000000";
      when "000111011011101" => color_data <= "000000000000";
      when "000111011011110" => color_data <= "000000000000";
      when "000111011011111" => color_data <= "000000000000";
      when "000111011100000" => color_data <= "000000000000";
      when "000111011100001" => color_data <= "000000000000";
      when "000111011100010" => color_data <= "000000000000";
      when "000111011100011" => color_data <= "000000000000";
      when "000111100000000" => color_data <= "000000000000";
      when "000111100000001" => color_data <= "000000000000";
      when "000111100000010" => color_data <= "000000000000";
      when "000111100000011" => color_data <= "000000000000";
      when "000111100000100" => color_data <= "000000000000";
      when "000111100000101" => color_data <= "000000000000";
      when "000111100000110" => color_data <= "000000000000";
      when "000111100000111" => color_data <= "000000000000";
      when "000111100001000" => color_data <= "000100010001";
      when "000111100001001" => color_data <= "001100100010";
      when "000111100001010" => color_data <= "001000100001";
      when "000111100001011" => color_data <= "001100110010";
      when "000111100001100" => color_data <= "001100110010";
      when "000111100001101" => color_data <= "001100110010";
      when "000111100001110" => color_data <= "001100110010";
      when "000111100001111" => color_data <= "001000100010";
      when "000111100010000" => color_data <= "001100100010";
      when "000111100010001" => color_data <= "000000000000";
      when "000111100010010" => color_data <= "000000000000";
      when "000111100010011" => color_data <= "000000000000";
      when "000111100010100" => color_data <= "000000000000";
      when "000111100010101" => color_data <= "100110000010";
      when "000111100010110" => color_data <= "111111000000";
      when "000111100010111" => color_data <= "111111010000";
      when "000111100011000" => color_data <= "111111010000";
      when "000111100011001" => color_data <= "111111010000";
      when "000111100011010" => color_data <= "111111010000";
      when "000111100011011" => color_data <= "111111010010";
      when "000111100011100" => color_data <= "111111111101";
      when "000111100011101" => color_data <= "111111111101";
      when "000111100011110" => color_data <= "111111111101";
      when "000111100011111" => color_data <= "111111111101";
      when "000111100100000" => color_data <= "111111111100";
      when "000111100100001" => color_data <= "111111111101";
      when "000111100100010" => color_data <= "111111111101";
      when "000111100100011" => color_data <= "111111111101";
      when "000111100100100" => color_data <= "111111111101";
      when "000111100100101" => color_data <= "111111111101";
      when "000111100100110" => color_data <= "111111111101";
      when "000111100100111" => color_data <= "111111111101";
      when "000111100101000" => color_data <= "111111111101";
      when "000111100101001" => color_data <= "111111111101";
      when "000111100101010" => color_data <= "111111111101";
      when "000111100101011" => color_data <= "111111111101";
      when "000111100101100" => color_data <= "111111111101";
      when "000111100101101" => color_data <= "111111111101";
      when "000111100101110" => color_data <= "111111111101";
      when "000111100101111" => color_data <= "111111111101";
      when "000111100110000" => color_data <= "111111111101";
      when "000111100110001" => color_data <= "111111111110";
      when "000111100110010" => color_data <= "111111111001";
      when "000111100110011" => color_data <= "111111100110";
      when "000111100110100" => color_data <= "111111100111";
      when "000111100110101" => color_data <= "111111100110";
      when "000111100110110" => color_data <= "111111100111";
      when "000111100110111" => color_data <= "111111100111";
      when "000111100111000" => color_data <= "111111100111";
      when "000111100111001" => color_data <= "111111100111";
      when "000111100111010" => color_data <= "111111100111";
      when "000111100111011" => color_data <= "111111100111";
      when "000111100111100" => color_data <= "111111100111";
      when "000111100111101" => color_data <= "111111100111";
      when "000111100111110" => color_data <= "111111100111";
      when "000111100111111" => color_data <= "111111100111";
      when "000111101000000" => color_data <= "111111100111";
      when "000111101000001" => color_data <= "111111100111";
      when "000111101000010" => color_data <= "111111100111";
      when "000111101000011" => color_data <= "111111100111";
      when "000111101000100" => color_data <= "111111100111";
      when "000111101000101" => color_data <= "111111100110";
      when "000111101000110" => color_data <= "111111100110";
      when "000111101000111" => color_data <= "111111100110";
      when "000111101001000" => color_data <= "111111100111";
      when "000111101001001" => color_data <= "111111100111";
      when "000111101001010" => color_data <= "111111010010";
      when "000111101001011" => color_data <= "111111010000";
      when "000111101001100" => color_data <= "111111010000";
      when "000111101001101" => color_data <= "111111010000";
      when "000111101001110" => color_data <= "111111000000";
      when "000111101001111" => color_data <= "011001100011";
      when "000111101010000" => color_data <= "000000000000";
      when "000111101010001" => color_data <= "000000000000";
      when "000111101010010" => color_data <= "000000000000";
      when "000111101010011" => color_data <= "000000000000";
      when "000111101010100" => color_data <= "000000000000";
      when "000111101010101" => color_data <= "000000000000";
      when "000111101010110" => color_data <= "000000000000";
      when "000111101010111" => color_data <= "000000000000";
      when "000111101011000" => color_data <= "000000000000";
      when "000111101011001" => color_data <= "000000000000";
      when "000111101011010" => color_data <= "000000000000";
      when "000111101011011" => color_data <= "000000000000";
      when "000111101011100" => color_data <= "000000000000";
      when "000111101011101" => color_data <= "000000000000";
      when "000111101011110" => color_data <= "000000000000";
      when "000111101011111" => color_data <= "000000000000";
      when "000111101100000" => color_data <= "000000000000";
      when "000111101100001" => color_data <= "000000000000";
      when "000111101100010" => color_data <= "000000000000";
      when "000111101100011" => color_data <= "000000000000";
      when "000111110000000" => color_data <= "000000000000";
      when "000111110000001" => color_data <= "000000000000";
      when "000111110000010" => color_data <= "000000000000";
      when "000111110000011" => color_data <= "000000000000";
      when "000111110000100" => color_data <= "000000000000";
      when "000111110000101" => color_data <= "000000000000";
      when "000111110000110" => color_data <= "000000000000";
      when "000111110000111" => color_data <= "000000000000";
      when "000111110001000" => color_data <= "110110100000";
      when "000111110001001" => color_data <= "111110110000";
      when "000111110001010" => color_data <= "111111000000";
      when "000111110001011" => color_data <= "110010100000";
      when "000111110001100" => color_data <= "110010100000";
      when "000111110001101" => color_data <= "110010100000";
      when "000111110001110" => color_data <= "110010010001";
      when "000111110001111" => color_data <= "110110100000";
      when "000111110010000" => color_data <= "111110110000";
      when "000111110010001" => color_data <= "010000110010";
      when "000111110010010" => color_data <= "000000000000";
      when "000111110010011" => color_data <= "000000000000";
      when "000111110010100" => color_data <= "000000000000";
      when "000111110010101" => color_data <= "110110110000";
      when "000111110010110" => color_data <= "111111010000";
      when "000111110010111" => color_data <= "111111010000";
      when "000111110011000" => color_data <= "111111010000";
      when "000111110011001" => color_data <= "111111010000";
      when "000111110011010" => color_data <= "111111010000";
      when "000111110011011" => color_data <= "111111010010";
      when "000111110011100" => color_data <= "111111111101";
      when "000111110011101" => color_data <= "111111111101";
      when "000111110011110" => color_data <= "111111111101";
      when "000111110011111" => color_data <= "111111111101";
      when "000111110100000" => color_data <= "111111111101";
      when "000111110100001" => color_data <= "111111111101";
      when "000111110100010" => color_data <= "111111111101";
      when "000111110100011" => color_data <= "111111111101";
      when "000111110100100" => color_data <= "111111111101";
      when "000111110100101" => color_data <= "111111111101";
      when "000111110100110" => color_data <= "111111111101";
      when "000111110100111" => color_data <= "111111111101";
      when "000111110101000" => color_data <= "111111111101";
      when "000111110101001" => color_data <= "111111111101";
      when "000111110101010" => color_data <= "111111111101";
      when "000111110101011" => color_data <= "111111111101";
      when "000111110101100" => color_data <= "111111111101";
      when "000111110101101" => color_data <= "111111111101";
      when "000111110101110" => color_data <= "111111111101";
      when "000111110101111" => color_data <= "111111111101";
      when "000111110110000" => color_data <= "111111111111";
      when "000111110110001" => color_data <= "111111111110";
      when "000111110110010" => color_data <= "111111100100";
      when "000111110110011" => color_data <= "111111010010";
      when "000111110110100" => color_data <= "111111100111";
      when "000111110110101" => color_data <= "111111100111";
      when "000111110110110" => color_data <= "111111100110";
      when "000111110110111" => color_data <= "111111100111";
      when "000111110111000" => color_data <= "111111100111";
      when "000111110111001" => color_data <= "111111100111";
      when "000111110111010" => color_data <= "111111100111";
      when "000111110111011" => color_data <= "111111100111";
      when "000111110111100" => color_data <= "111111100111";
      when "000111110111101" => color_data <= "111111100111";
      when "000111110111110" => color_data <= "111111100111";
      when "000111110111111" => color_data <= "111111100111";
      when "000111111000000" => color_data <= "111111100111";
      when "000111111000001" => color_data <= "111111100111";
      when "000111111000010" => color_data <= "111111100111";
      when "000111111000011" => color_data <= "111111100111";
      when "000111111000100" => color_data <= "111111100111";
      when "000111111000101" => color_data <= "111111100111";
      when "000111111000110" => color_data <= "111111100111";
      when "000111111000111" => color_data <= "111111100111";
      when "000111111001000" => color_data <= "111111100111";
      when "000111111001001" => color_data <= "111111100111";
      when "000111111001010" => color_data <= "111111010011";
      when "000111111001011" => color_data <= "111111010000";
      when "000111111001100" => color_data <= "111111010000";
      when "000111111001101" => color_data <= "111111010000";
      when "000111111001110" => color_data <= "111111000000";
      when "000111111001111" => color_data <= "101010000010";
      when "000111111010000" => color_data <= "000000000000";
      when "000111111010001" => color_data <= "000000000000";
      when "000111111010010" => color_data <= "000000000000";
      when "000111111010011" => color_data <= "000000000000";
      when "000111111010100" => color_data <= "000000000000";
      when "000111111010101" => color_data <= "000000000000";
      when "000111111010110" => color_data <= "100001110010";
      when "000111111010111" => color_data <= "100001100010";
      when "000111111011000" => color_data <= "100101110010";
      when "000111111011001" => color_data <= "100110000010";
      when "000111111011010" => color_data <= "100110000010";
      when "000111111011011" => color_data <= "100110000010";
      when "000111111011100" => color_data <= "011101100011";
      when "000111111011101" => color_data <= "011101100011";
      when "000111111011110" => color_data <= "011101100011";
      when "000111111011111" => color_data <= "000000000000";
      when "000111111100000" => color_data <= "000000000000";
      when "000111111100001" => color_data <= "000000000000";
      when "000111111100010" => color_data <= "000000000000";
      when "000111111100011" => color_data <= "000000000000";
      when "001000000000000" => color_data <= "000000000000";
      when "001000000000001" => color_data <= "000000000000";
      when "001000000000010" => color_data <= "000000000000";
      when "001000000000011" => color_data <= "000000000000";
      when "001000000000100" => color_data <= "000000000000";
      when "001000000000101" => color_data <= "000000000000";
      when "001000000000110" => color_data <= "000000000000";
      when "001000000000111" => color_data <= "001100110010";
      when "001000000001000" => color_data <= "111110110000";
      when "001000000001001" => color_data <= "111111000000";
      when "001000000001010" => color_data <= "111111000000";
      when "001000000001011" => color_data <= "001000100001";
      when "001000000001100" => color_data <= "000000000000";
      when "001000000001101" => color_data <= "000000000000";
      when "001000000001110" => color_data <= "000000000000";
      when "001000000001111" => color_data <= "101110010001";
      when "001000000010000" => color_data <= "111110110000";
      when "001000000010001" => color_data <= "001000010001";
      when "001000000010010" => color_data <= "000000000000";
      when "001000000010011" => color_data <= "000000000000";
      when "001000000010100" => color_data <= "001100110010";
      when "001000000010101" => color_data <= "111111000000";
      when "001000000010110" => color_data <= "111111010000";
      when "001000000010111" => color_data <= "111111010000";
      when "001000000011000" => color_data <= "111111010000";
      when "001000000011001" => color_data <= "111111010000";
      when "001000000011010" => color_data <= "111111010000";
      when "001000000011011" => color_data <= "111111010010";
      when "001000000011100" => color_data <= "111111111101";
      when "001000000011101" => color_data <= "111111111101";
      when "001000000011110" => color_data <= "111111111101";
      when "001000000011111" => color_data <= "111111111101";
      when "001000000100000" => color_data <= "111111111101";
      when "001000000100001" => color_data <= "111111111101";
      when "001000000100010" => color_data <= "111111111101";
      when "001000000100011" => color_data <= "111111111101";
      when "001000000100100" => color_data <= "111111111101";
      when "001000000100101" => color_data <= "111111111101";
      when "001000000100110" => color_data <= "111111111101";
      when "001000000100111" => color_data <= "111111111101";
      when "001000000101000" => color_data <= "111111111101";
      when "001000000101001" => color_data <= "111111111101";
      when "001000000101010" => color_data <= "111111111101";
      when "001000000101011" => color_data <= "111111111101";
      when "001000000101100" => color_data <= "111111111101";
      when "001000000101101" => color_data <= "111111111100";
      when "001000000101110" => color_data <= "111111111101";
      when "001000000101111" => color_data <= "111111111111";
      when "001000000110000" => color_data <= "111111111011";
      when "001000000110001" => color_data <= "111111010010";
      when "001000000110010" => color_data <= "111111000000";
      when "001000000110011" => color_data <= "111111010000";
      when "001000000110100" => color_data <= "111111010001";
      when "001000000110101" => color_data <= "111111100110";
      when "001000000110110" => color_data <= "111111101000";
      when "001000000110111" => color_data <= "111111100111";
      when "001000000111000" => color_data <= "111111100110";
      when "001000000111001" => color_data <= "111111100111";
      when "001000000111010" => color_data <= "111111100111";
      when "001000000111011" => color_data <= "111111100111";
      when "001000000111100" => color_data <= "111111100111";
      when "001000000111101" => color_data <= "111111100111";
      when "001000000111110" => color_data <= "111111100111";
      when "001000000111111" => color_data <= "111111100111";
      when "001000001000000" => color_data <= "111111100111";
      when "001000001000001" => color_data <= "111111100111";
      when "001000001000010" => color_data <= "111111100111";
      when "001000001000011" => color_data <= "111111100111";
      when "001000001000100" => color_data <= "111111100111";
      when "001000001000101" => color_data <= "111111100111";
      when "001000001000110" => color_data <= "111111100111";
      when "001000001000111" => color_data <= "111111100111";
      when "001000001001000" => color_data <= "111111100111";
      when "001000001001001" => color_data <= "111111100111";
      when "001000001001010" => color_data <= "111111010010";
      when "001000001001011" => color_data <= "111111010000";
      when "001000001001100" => color_data <= "111111010000";
      when "001000001001101" => color_data <= "111111010000";
      when "001000001001110" => color_data <= "111111010000";
      when "001000001001111" => color_data <= "110010100000";
      when "001000001010000" => color_data <= "000000000000";
      when "001000001010001" => color_data <= "000000000000";
      when "001000001010010" => color_data <= "000000000000";
      when "001000001010011" => color_data <= "000000000000";
      when "001000001010100" => color_data <= "000000000000";
      when "001000001010101" => color_data <= "000000000000";
      when "001000001010110" => color_data <= "110110100000";
      when "001000001010111" => color_data <= "111110110000";
      when "001000001011000" => color_data <= "100001110010";
      when "001000001011001" => color_data <= "011101100011";
      when "001000001011010" => color_data <= "011101100010";
      when "001000001011011" => color_data <= "100001110010";
      when "001000001011100" => color_data <= "110110100000";
      when "001000001011101" => color_data <= "111110110000";
      when "001000001011110" => color_data <= "111110110000";
      when "001000001011111" => color_data <= "010101010011";
      when "001000001100000" => color_data <= "000000000000";
      when "001000001100001" => color_data <= "000000000000";
      when "001000001100010" => color_data <= "000000000000";
      when "001000001100011" => color_data <= "000000000000";
      when "001000010000000" => color_data <= "000000000000";
      when "001000010000001" => color_data <= "000000000000";
      when "001000010000010" => color_data <= "000000000000";
      when "001000010000011" => color_data <= "000000000000";
      when "001000010000100" => color_data <= "000000000000";
      when "001000010000101" => color_data <= "000000000000";
      when "001000010000110" => color_data <= "000000000000";
      when "001000010000111" => color_data <= "001100110010";
      when "001000010001000" => color_data <= "111110110000";
      when "001000010001001" => color_data <= "111111000000";
      when "001000010001010" => color_data <= "111111000000";
      when "001000010001011" => color_data <= "000000000000";
      when "001000010001100" => color_data <= "000000000000";
      when "001000010001101" => color_data <= "000000000000";
      when "001000010001110" => color_data <= "000100010001";
      when "001000010001111" => color_data <= "110110100000";
      when "001000010010000" => color_data <= "111110110000";
      when "001000010010001" => color_data <= "001000100001";
      when "001000010010010" => color_data <= "000000000000";
      when "001000010010011" => color_data <= "000000000000";
      when "001000010010100" => color_data <= "010101010011";
      when "001000010010101" => color_data <= "111111000000";
      when "001000010010110" => color_data <= "111111010000";
      when "001000010010111" => color_data <= "111111010000";
      when "001000010011000" => color_data <= "111111010000";
      when "001000010011001" => color_data <= "111111010000";
      when "001000010011010" => color_data <= "111111010000";
      when "001000010011011" => color_data <= "111111010010";
      when "001000010011100" => color_data <= "111111111101";
      when "001000010011101" => color_data <= "111111111110";
      when "001000010011110" => color_data <= "111111111100";
      when "001000010011111" => color_data <= "111111111101";
      when "001000010100000" => color_data <= "111111111101";
      when "001000010100001" => color_data <= "111111111101";
      when "001000010100010" => color_data <= "111111111101";
      when "001000010100011" => color_data <= "111111111101";
      when "001000010100100" => color_data <= "111111111101";
      when "001000010100101" => color_data <= "111111111101";
      when "001000010100110" => color_data <= "111111111101";
      when "001000010100111" => color_data <= "111111111101";
      when "001000010101000" => color_data <= "111111111101";
      when "001000010101001" => color_data <= "111111111101";
      when "001000010101010" => color_data <= "111111111101";
      when "001000010101011" => color_data <= "111111111101";
      when "001000010101100" => color_data <= "111111111101";
      when "001000010101101" => color_data <= "111111111110";
      when "001000010101110" => color_data <= "111111111110";
      when "001000010101111" => color_data <= "111111100111";
      when "001000010110000" => color_data <= "111111010000";
      when "001000010110001" => color_data <= "111111000000";
      when "001000010110010" => color_data <= "111111010000";
      when "001000010110011" => color_data <= "111111010001";
      when "001000010110100" => color_data <= "111111010000";
      when "001000010110101" => color_data <= "111111010000";
      when "001000010110110" => color_data <= "111111010100";
      when "001000010110111" => color_data <= "111111101000";
      when "001000010111000" => color_data <= "111111100111";
      when "001000010111001" => color_data <= "111111100111";
      when "001000010111010" => color_data <= "111111100111";
      when "001000010111011" => color_data <= "111111100111";
      when "001000010111100" => color_data <= "111111100111";
      when "001000010111101" => color_data <= "111111100111";
      when "001000010111110" => color_data <= "111111100111";
      when "001000010111111" => color_data <= "111111100111";
      when "001000011000000" => color_data <= "111111100111";
      when "001000011000001" => color_data <= "111111100111";
      when "001000011000010" => color_data <= "111111100111";
      when "001000011000011" => color_data <= "111111100111";
      when "001000011000100" => color_data <= "111111100111";
      when "001000011000101" => color_data <= "111111100111";
      when "001000011000110" => color_data <= "111111100111";
      when "001000011000111" => color_data <= "111111100111";
      when "001000011001000" => color_data <= "111111100111";
      when "001000011001001" => color_data <= "111111100111";
      when "001000011001010" => color_data <= "111111010010";
      when "001000011001011" => color_data <= "111111010000";
      when "001000011001100" => color_data <= "111111010000";
      when "001000011001101" => color_data <= "111111010000";
      when "001000011001110" => color_data <= "111111010000";
      when "001000011001111" => color_data <= "110110110000";
      when "001000011010000" => color_data <= "001000100001";
      when "001000011010001" => color_data <= "000000000000";
      when "001000011010010" => color_data <= "000000000000";
      when "001000011010011" => color_data <= "000000000000";
      when "001000011010100" => color_data <= "000000000000";
      when "001000011010101" => color_data <= "000000000000";
      when "001000011010110" => color_data <= "110010010001";
      when "001000011010111" => color_data <= "111110110000";
      when "001000011011000" => color_data <= "000100010000";
      when "001000011011001" => color_data <= "000000000000";
      when "001000011011010" => color_data <= "000000000000";
      when "001000011011011" => color_data <= "000000000000";
      when "001000011011100" => color_data <= "101110010001";
      when "001000011011101" => color_data <= "111111000000";
      when "001000011011110" => color_data <= "111110110000";
      when "001000011011111" => color_data <= "011001010011";
      when "001000011100000" => color_data <= "000000000000";
      when "001000011100001" => color_data <= "000000000000";
      when "001000011100010" => color_data <= "000000000000";
      when "001000011100011" => color_data <= "000000000000";
      when "001000100000000" => color_data <= "000000000000";
      when "001000100000001" => color_data <= "000000000000";
      when "001000100000010" => color_data <= "000000000000";
      when "001000100000011" => color_data <= "000000000000";
      when "001000100000100" => color_data <= "000000000000";
      when "001000100000101" => color_data <= "000000000000";
      when "001000100000110" => color_data <= "000000000000";
      when "001000100000111" => color_data <= "001100100010";
      when "001000100001000" => color_data <= "111110110000";
      when "001000100001001" => color_data <= "111111000000";
      when "001000100001010" => color_data <= "111111000000";
      when "001000100001011" => color_data <= "000000000000";
      when "001000100001100" => color_data <= "000000000000";
      when "001000100001101" => color_data <= "000000000000";
      when "001000100001110" => color_data <= "000100010001";
      when "001000100001111" => color_data <= "110110100000";
      when "001000100010000" => color_data <= "111110110000";
      when "001000100010001" => color_data <= "011101100011";
      when "001000100010010" => color_data <= "000000000000";
      when "001000100010011" => color_data <= "000000000000";
      when "001000100010100" => color_data <= "100001110010";
      when "001000100010101" => color_data <= "111111000000";
      when "001000100010110" => color_data <= "111111010000";
      when "001000100010111" => color_data <= "111111010000";
      when "001000100011000" => color_data <= "111111010000";
      when "001000100011001" => color_data <= "111111010000";
      when "001000100011010" => color_data <= "111111010000";
      when "001000100011011" => color_data <= "111111010000";
      when "001000100011100" => color_data <= "111111111001";
      when "001000100011101" => color_data <= "111111111110";
      when "001000100011110" => color_data <= "111111111110";
      when "001000100011111" => color_data <= "111111111101";
      when "001000100100000" => color_data <= "111111111101";
      when "001000100100001" => color_data <= "111111111101";
      when "001000100100010" => color_data <= "111111111101";
      when "001000100100011" => color_data <= "111111111101";
      when "001000100100100" => color_data <= "111111111101";
      when "001000100100101" => color_data <= "111111111101";
      when "001000100100110" => color_data <= "111111111101";
      when "001000100100111" => color_data <= "111111111101";
      when "001000100101000" => color_data <= "111111111101";
      when "001000100101001" => color_data <= "111111111101";
      when "001000100101010" => color_data <= "111111111100";
      when "001000100101011" => color_data <= "111111111101";
      when "001000100101100" => color_data <= "111111111111";
      when "001000100101101" => color_data <= "111111111011";
      when "001000100101110" => color_data <= "111111010010";
      when "001000100101111" => color_data <= "111111000000";
      when "001000100110000" => color_data <= "111111010000";
      when "001000100110001" => color_data <= "111111010001";
      when "001000100110010" => color_data <= "111111010000";
      when "001000100110011" => color_data <= "111111010000";
      when "001000100110100" => color_data <= "111111010001";
      when "001000100110101" => color_data <= "111111010000";
      when "001000100110110" => color_data <= "111111010000";
      when "001000100110111" => color_data <= "111111010010";
      when "001000100111000" => color_data <= "111111100111";
      when "001000100111001" => color_data <= "111111101000";
      when "001000100111010" => color_data <= "111111100111";
      when "001000100111011" => color_data <= "111111100111";
      when "001000100111100" => color_data <= "111111100111";
      when "001000100111101" => color_data <= "111111100111";
      when "001000100111110" => color_data <= "111111100111";
      when "001000100111111" => color_data <= "111111100111";
      when "001000101000000" => color_data <= "111111100111";
      when "001000101000001" => color_data <= "111111100111";
      when "001000101000010" => color_data <= "111111100111";
      when "001000101000011" => color_data <= "111111100111";
      when "001000101000100" => color_data <= "111111100111";
      when "001000101000101" => color_data <= "111111100111";
      when "001000101000110" => color_data <= "111111100111";
      when "001000101000111" => color_data <= "111111100111";
      when "001000101001000" => color_data <= "111111100111";
      when "001000101001001" => color_data <= "111111100111";
      when "001000101001010" => color_data <= "111111010001";
      when "001000101001011" => color_data <= "111111010000";
      when "001000101001100" => color_data <= "111111010000";
      when "001000101001101" => color_data <= "111111010000";
      when "001000101001110" => color_data <= "111111010000";
      when "001000101001111" => color_data <= "111111000000";
      when "001000101010000" => color_data <= "010101010011";
      when "001000101010001" => color_data <= "000000000000";
      when "001000101010010" => color_data <= "000000000000";
      when "001000101010011" => color_data <= "000000000000";
      when "001000101010100" => color_data <= "000000000000";
      when "001000101010101" => color_data <= "000100010001";
      when "001000101010110" => color_data <= "110110100000";
      when "001000101010111" => color_data <= "111110110000";
      when "001000101011000" => color_data <= "010101000010";
      when "001000101011001" => color_data <= "000000000000";
      when "001000101011010" => color_data <= "000000000000";
      when "001000101011011" => color_data <= "000000000000";
      when "001000101011100" => color_data <= "101010000010";
      when "001000101011101" => color_data <= "111111000000";
      when "001000101011110" => color_data <= "111110110000";
      when "001000101011111" => color_data <= "011001010011";
      when "001000101100000" => color_data <= "000000000000";
      when "001000101100001" => color_data <= "000000000000";
      when "001000101100010" => color_data <= "000000000000";
      when "001000101100011" => color_data <= "000000000000";
      when "001000110000000" => color_data <= "000000000000";
      when "001000110000001" => color_data <= "000000000000";
      when "001000110000010" => color_data <= "000000000000";
      when "001000110000011" => color_data <= "000000000000";
      when "001000110000100" => color_data <= "000000000000";
      when "001000110000101" => color_data <= "000000000000";
      when "001000110000110" => color_data <= "000000000000";
      when "001000110000111" => color_data <= "001000100001";
      when "001000110001000" => color_data <= "111111000000";
      when "001000110001001" => color_data <= "111111000000";
      when "001000110001010" => color_data <= "111111000000";
      when "001000110001011" => color_data <= "000100010001";
      when "001000110001100" => color_data <= "000000000000";
      when "001000110001101" => color_data <= "000000000000";
      when "001000110001110" => color_data <= "000000000000";
      when "001000110001111" => color_data <= "101010000010";
      when "001000110010000" => color_data <= "111110110000";
      when "001000110010001" => color_data <= "110110100000";
      when "001000110010010" => color_data <= "000100010001";
      when "001000110010011" => color_data <= "000000000000";
      when "001000110010100" => color_data <= "101010010010";
      when "001000110010101" => color_data <= "111111010000";
      when "001000110010110" => color_data <= "111111010001";
      when "001000110010111" => color_data <= "111111010000";
      when "001000110011000" => color_data <= "111111010000";
      when "001000110011001" => color_data <= "111111010000";
      when "001000110011010" => color_data <= "111111010000";
      when "001000110011011" => color_data <= "111111100101";
      when "001000110011100" => color_data <= "111111101000";
      when "001000110011101" => color_data <= "111111100111";
      when "001000110011110" => color_data <= "111111101010";
      when "001000110011111" => color_data <= "111111111100";
      when "001000110100000" => color_data <= "111111111110";
      when "001000110100001" => color_data <= "111111111101";
      when "001000110100010" => color_data <= "111111111101";
      when "001000110100011" => color_data <= "111111111101";
      when "001000110100100" => color_data <= "111111111101";
      when "001000110100101" => color_data <= "111111111101";
      when "001000110100110" => color_data <= "111111111101";
      when "001000110100111" => color_data <= "111111111101";
      when "001000110101000" => color_data <= "111111111100";
      when "001000110101001" => color_data <= "111111111101";
      when "001000110101010" => color_data <= "111111111111";
      when "001000110101011" => color_data <= "111111111110";
      when "001000110101100" => color_data <= "111111100111";
      when "001000110101101" => color_data <= "111111000000";
      when "001000110101110" => color_data <= "111111000000";
      when "001000110101111" => color_data <= "111111010000";
      when "001000110110000" => color_data <= "111111010001";
      when "001000110110001" => color_data <= "111111010000";
      when "001000110110010" => color_data <= "111111010000";
      when "001000110110011" => color_data <= "111111010000";
      when "001000110110100" => color_data <= "111111010000";
      when "001000110110101" => color_data <= "111111010000";
      when "001000110110110" => color_data <= "111111010000";
      when "001000110110111" => color_data <= "111111010000";
      when "001000110111000" => color_data <= "111111010001";
      when "001000110111001" => color_data <= "111111100101";
      when "001000110111010" => color_data <= "111111101000";
      when "001000110111011" => color_data <= "111111100111";
      when "001000110111100" => color_data <= "111111100110";
      when "001000110111101" => color_data <= "111111100111";
      when "001000110111110" => color_data <= "111111100111";
      when "001000110111111" => color_data <= "111111100111";
      when "001000111000000" => color_data <= "111111100111";
      when "001000111000001" => color_data <= "111111100111";
      when "001000111000010" => color_data <= "111111100111";
      when "001000111000011" => color_data <= "111111100111";
      when "001000111000100" => color_data <= "111111100111";
      when "001000111000101" => color_data <= "111111100111";
      when "001000111000110" => color_data <= "111111100111";
      when "001000111000111" => color_data <= "111111100111";
      when "001000111001000" => color_data <= "111111100111";
      when "001000111001001" => color_data <= "111111010101";
      when "001000111001010" => color_data <= "111111010000";
      when "001000111001011" => color_data <= "111111010000";
      when "001000111001100" => color_data <= "111111010000";
      when "001000111001101" => color_data <= "111111010000";
      when "001000111001110" => color_data <= "111111010000";
      when "001000111001111" => color_data <= "111111000000";
      when "001000111010000" => color_data <= "011101100011";
      when "001000111010001" => color_data <= "000000000000";
      when "001000111010010" => color_data <= "000000000000";
      when "001000111010011" => color_data <= "000000000000";
      when "001000111010100" => color_data <= "000000000000";
      when "001000111010101" => color_data <= "011101100011";
      when "001000111010110" => color_data <= "111110110000";
      when "001000111010111" => color_data <= "110110100000";
      when "001000111011000" => color_data <= "001000100010";
      when "001000111011001" => color_data <= "000000000000";
      when "001000111011010" => color_data <= "000000000000";
      when "001000111011011" => color_data <= "000000000000";
      when "001000111011100" => color_data <= "101110000001";
      when "001000111011101" => color_data <= "111111000000";
      when "001000111011110" => color_data <= "111110110000";
      when "001000111011111" => color_data <= "010101010010";
      when "001000111100000" => color_data <= "000000000000";
      when "001000111100001" => color_data <= "000000000000";
      when "001000111100010" => color_data <= "000000000000";
      when "001000111100011" => color_data <= "000000000000";
      when "001001000000000" => color_data <= "000000000000";
      when "001001000000001" => color_data <= "000000000000";
      when "001001000000010" => color_data <= "000000000000";
      when "001001000000011" => color_data <= "000000000000";
      when "001001000000100" => color_data <= "000000000000";
      when "001001000000101" => color_data <= "000000000000";
      when "001001000000110" => color_data <= "000000000000";
      when "001001000000111" => color_data <= "000100010001";
      when "001001000001000" => color_data <= "110110100000";
      when "001001000001001" => color_data <= "111111000000";
      when "001001000001010" => color_data <= "111110110000";
      when "001001000001011" => color_data <= "001000100010";
      when "001001000001100" => color_data <= "000000000000";
      when "001001000001101" => color_data <= "000000000000";
      when "001001000001110" => color_data <= "000000000000";
      when "001001000001111" => color_data <= "010001000010";
      when "001001000010000" => color_data <= "110110100000";
      when "001001000010001" => color_data <= "111111000000";
      when "001001000010010" => color_data <= "110010010000";
      when "001001000010011" => color_data <= "001100110010";
      when "001001000010100" => color_data <= "101010010010";
      when "001001000010101" => color_data <= "111111010000";
      when "001001000010110" => color_data <= "111111010000";
      when "001001000010111" => color_data <= "111111010000";
      when "001001000011000" => color_data <= "111111010000";
      when "001001000011001" => color_data <= "111111010000";
      when "001001000011010" => color_data <= "111111100100";
      when "001001000011011" => color_data <= "111111111011";
      when "001001000011100" => color_data <= "111111111011";
      when "001001000011101" => color_data <= "111111101000";
      when "001001000011110" => color_data <= "111111100111";
      when "001001000011111" => color_data <= "111111100111";
      when "001001000100000" => color_data <= "111111101001";
      when "001001000100001" => color_data <= "111111111010";
      when "001001000100010" => color_data <= "111111111100";
      when "001001000100011" => color_data <= "111111111110";
      when "001001000100100" => color_data <= "111111111110";
      when "001001000100101" => color_data <= "111111111101";
      when "001001000100110" => color_data <= "111111111101";
      when "001001000100111" => color_data <= "111111111100";
      when "001001000101000" => color_data <= "111111111101";
      when "001001000101001" => color_data <= "111111111111";
      when "001001000101010" => color_data <= "111111111011";
      when "001001000101011" => color_data <= "111111010010";
      when "001001000101100" => color_data <= "111111000000";
      when "001001000101101" => color_data <= "111111010000";
      when "001001000101110" => color_data <= "111111010001";
      when "001001000101111" => color_data <= "111111010000";
      when "001001000110000" => color_data <= "111111010000";
      when "001001000110001" => color_data <= "111111010000";
      when "001001000110010" => color_data <= "111111010000";
      when "001001000110011" => color_data <= "111111010000";
      when "001001000110100" => color_data <= "111111010000";
      when "001001000110101" => color_data <= "111111010000";
      when "001001000110110" => color_data <= "111111010000";
      when "001001000110111" => color_data <= "111111010000";
      when "001001000111000" => color_data <= "111111010000";
      when "001001000111001" => color_data <= "111111010000";
      when "001001000111010" => color_data <= "111111010011";
      when "001001000111011" => color_data <= "111111100111";
      when "001001000111100" => color_data <= "111111100111";
      when "001001000111101" => color_data <= "111111100111";
      when "001001000111110" => color_data <= "111111100111";
      when "001001000111111" => color_data <= "111111100111";
      when "001001001000000" => color_data <= "111111100111";
      when "001001001000001" => color_data <= "111111100111";
      when "001001001000010" => color_data <= "111111100111";
      when "001001001000011" => color_data <= "111111100111";
      when "001001001000100" => color_data <= "111111100111";
      when "001001001000101" => color_data <= "111111100111";
      when "001001001000110" => color_data <= "111111100111";
      when "001001001000111" => color_data <= "111111100101";
      when "001001001001000" => color_data <= "111111100100";
      when "001001001001001" => color_data <= "111111100111";
      when "001001001001010" => color_data <= "111111010011";
      when "001001001001011" => color_data <= "111111010000";
      when "001001001001100" => color_data <= "111111010000";
      when "001001001001101" => color_data <= "111111010000";
      when "001001001001110" => color_data <= "111111010000";
      when "001001001001111" => color_data <= "111111000000";
      when "001001001010000" => color_data <= "100001110010";
      when "001001001010001" => color_data <= "000000000000";
      when "001001001010010" => color_data <= "000000000000";
      when "001001001010011" => color_data <= "000000000000";
      when "001001001010100" => color_data <= "010001000010";
      when "001001001010101" => color_data <= "110110100000";
      when "001001001010110" => color_data <= "111110110000";
      when "001001001010111" => color_data <= "101110010001";
      when "001001001011000" => color_data <= "000000000000";
      when "001001001011001" => color_data <= "000000000000";
      when "001001001011010" => color_data <= "000000000000";
      when "001001001011011" => color_data <= "000000000000";
      when "001001001011100" => color_data <= "110010010001";
      when "001001001011101" => color_data <= "111111000000";
      when "001001001011110" => color_data <= "111110110000";
      when "001001001011111" => color_data <= "010001000010";
      when "001001001100000" => color_data <= "000000000000";
      when "001001001100001" => color_data <= "000000000000";
      when "001001001100010" => color_data <= "000000000000";
      when "001001001100011" => color_data <= "000000000000";
      when "001001010000000" => color_data <= "000000000000";
      when "001001010000001" => color_data <= "000000000000";
      when "001001010000010" => color_data <= "000000000000";
      when "001001010000011" => color_data <= "000000000000";
      when "001001010000100" => color_data <= "000000000000";
      when "001001010000101" => color_data <= "000000000000";
      when "001001010000110" => color_data <= "000000000000";
      when "001001010000111" => color_data <= "000000000000";
      when "001001010001000" => color_data <= "110010010001";
      when "001001010001001" => color_data <= "111111000000";
      when "001001010001010" => color_data <= "111110110000";
      when "001001010001011" => color_data <= "010001000010";
      when "001001010001100" => color_data <= "000000000000";
      when "001001010001101" => color_data <= "000000000000";
      when "001001010001110" => color_data <= "000000000000";
      when "001001010001111" => color_data <= "000000000000";
      when "001001010010000" => color_data <= "101110010001";
      when "001001010010001" => color_data <= "111110110000";
      when "001001010010010" => color_data <= "111111000000";
      when "001001010010011" => color_data <= "111111000000";
      when "001001010010100" => color_data <= "111111010001";
      when "001001010010101" => color_data <= "111111010000";
      when "001001010010110" => color_data <= "111111010000";
      when "001001010010111" => color_data <= "111111010001";
      when "001001010011000" => color_data <= "111111000000";
      when "001001010011001" => color_data <= "111111010011";
      when "001001010011010" => color_data <= "111111111011";
      when "001001010011011" => color_data <= "111111101010";
      when "001001010011100" => color_data <= "111111101001";
      when "001001010011101" => color_data <= "111111101010";
      when "001001010011110" => color_data <= "111111101010";
      when "001001010011111" => color_data <= "111111101001";
      when "001001010100000" => color_data <= "111111100111";
      when "001001010100001" => color_data <= "111111100110";
      when "001001010100010" => color_data <= "111111101000";
      when "001001010100011" => color_data <= "111111101001";
      when "001001010100100" => color_data <= "111111111010";
      when "001001010100101" => color_data <= "111111111100";
      when "001001010100110" => color_data <= "111111111101";
      when "001001010100111" => color_data <= "111111111111";
      when "001001010101000" => color_data <= "111111111110";
      when "001001010101001" => color_data <= "111111100111";
      when "001001010101010" => color_data <= "111111000000";
      when "001001010101011" => color_data <= "111111000000";
      when "001001010101100" => color_data <= "111111010000";
      when "001001010101101" => color_data <= "111111010000";
      when "001001010101110" => color_data <= "111111010000";
      when "001001010101111" => color_data <= "111111010000";
      when "001001010110000" => color_data <= "111111010000";
      when "001001010110001" => color_data <= "111111010000";
      when "001001010110010" => color_data <= "111111010000";
      when "001001010110011" => color_data <= "111111010000";
      when "001001010110100" => color_data <= "111111010000";
      when "001001010110101" => color_data <= "111111010000";
      when "001001010110110" => color_data <= "111111010000";
      when "001001010110111" => color_data <= "111111010000";
      when "001001010111000" => color_data <= "111111010000";
      when "001001010111001" => color_data <= "111111010000";
      when "001001010111010" => color_data <= "111111010000";
      when "001001010111011" => color_data <= "111111010001";
      when "001001010111100" => color_data <= "111111100110";
      when "001001010111101" => color_data <= "111111101000";
      when "001001010111110" => color_data <= "111111100111";
      when "001001010111111" => color_data <= "111111100111";
      when "001001011000000" => color_data <= "111111100111";
      when "001001011000001" => color_data <= "111111100110";
      when "001001011000010" => color_data <= "111111100111";
      when "001001011000011" => color_data <= "111111100111";
      when "001001011000100" => color_data <= "111111100110";
      when "001001011000101" => color_data <= "111111100101";
      when "001001011000110" => color_data <= "111111010101";
      when "001001011000111" => color_data <= "111111100110";
      when "001001011001000" => color_data <= "111111101000";
      when "001001011001001" => color_data <= "111111111011";
      when "001001011001010" => color_data <= "111111101001";
      when "001001011001011" => color_data <= "111111010000";
      when "001001011001100" => color_data <= "111111010000";
      when "001001011001101" => color_data <= "111111010000";
      when "001001011001110" => color_data <= "111111010000";
      when "001001011001111" => color_data <= "111111000000";
      when "001001011010000" => color_data <= "100001110010";
      when "001001011010001" => color_data <= "000000000000";
      when "001001011010010" => color_data <= "000000000000";
      when "001001011010011" => color_data <= "010101010011";
      when "001001011010100" => color_data <= "110110100000";
      when "001001011010101" => color_data <= "111111000000";
      when "001001011010110" => color_data <= "110110100000";
      when "001001011010111" => color_data <= "010101000010";
      when "001001011011000" => color_data <= "000000000000";
      when "001001011011001" => color_data <= "000000000000";
      when "001001011011010" => color_data <= "000000000000";
      when "001001011011011" => color_data <= "000000000000";
      when "001001011011100" => color_data <= "110110100000";
      when "001001011011101" => color_data <= "111111000000";
      when "001001011011110" => color_data <= "111110110000";
      when "001001011011111" => color_data <= "001100110010";
      when "001001011100000" => color_data <= "000000000000";
      when "001001011100001" => color_data <= "000000000000";
      when "001001011100010" => color_data <= "000000000000";
      when "001001011100011" => color_data <= "000000000000";
      when "001001100000000" => color_data <= "000000000000";
      when "001001100000001" => color_data <= "000000000000";
      when "001001100000010" => color_data <= "000000000000";
      when "001001100000011" => color_data <= "000000000000";
      when "001001100000100" => color_data <= "000000000000";
      when "001001100000101" => color_data <= "000000000000";
      when "001001100000110" => color_data <= "000000000000";
      when "001001100000111" => color_data <= "000000000000";
      when "001001100001000" => color_data <= "100110000010";
      when "001001100001001" => color_data <= "111110110000";
      when "001001100001010" => color_data <= "111110110000";
      when "001001100001011" => color_data <= "011101100011";
      when "001001100001100" => color_data <= "000000000000";
      when "001001100001101" => color_data <= "000000000000";
      when "001001100001110" => color_data <= "000000000000";
      when "001001100001111" => color_data <= "000000000000";
      when "001001100010000" => color_data <= "000100010001";
      when "001001100010001" => color_data <= "110110100000";
      when "001001100010010" => color_data <= "111111000000";
      when "001001100010011" => color_data <= "111111000000";
      when "001001100010100" => color_data <= "111111010000";
      when "001001100010101" => color_data <= "111111010000";
      when "001001100010110" => color_data <= "111111010000";
      when "001001100010111" => color_data <= "111111000000";
      when "001001100011000" => color_data <= "111111010010";
      when "001001100011001" => color_data <= "111111111010";
      when "001001100011010" => color_data <= "111111101011";
      when "001001100011011" => color_data <= "111111101001";
      when "001001100011100" => color_data <= "111111101010";
      when "001001100011101" => color_data <= "111111101010";
      when "001001100011110" => color_data <= "111111101010";
      when "001001100011111" => color_data <= "111111101010";
      when "001001100100000" => color_data <= "111111101010";
      when "001001100100001" => color_data <= "111111101010";
      when "001001100100010" => color_data <= "111111101001";
      when "001001100100011" => color_data <= "111111100111";
      when "001001100100100" => color_data <= "111111100111";
      when "001001100100101" => color_data <= "111111101000";
      when "001001100100110" => color_data <= "111111101001";
      when "001001100100111" => color_data <= "111111111001";
      when "001001100101000" => color_data <= "111111010100";
      when "001001100101001" => color_data <= "111111000000";
      when "001001100101010" => color_data <= "111111010000";
      when "001001100101011" => color_data <= "111111010000";
      when "001001100101100" => color_data <= "111111010000";
      when "001001100101101" => color_data <= "111111010000";
      when "001001100101110" => color_data <= "111111010000";
      when "001001100101111" => color_data <= "111111010000";
      when "001001100110000" => color_data <= "111111010000";
      when "001001100110001" => color_data <= "111111010000";
      when "001001100110010" => color_data <= "111111010000";
      when "001001100110011" => color_data <= "111111010000";
      when "001001100110100" => color_data <= "111111010000";
      when "001001100110101" => color_data <= "111111010000";
      when "001001100110110" => color_data <= "111111010000";
      when "001001100110111" => color_data <= "111111010000";
      when "001001100111000" => color_data <= "111111010000";
      when "001001100111001" => color_data <= "111111010000";
      when "001001100111010" => color_data <= "111111010000";
      when "001001100111011" => color_data <= "111111010000";
      when "001001100111100" => color_data <= "111111010000";
      when "001001100111101" => color_data <= "111111010100";
      when "001001100111110" => color_data <= "111111101000";
      when "001001100111111" => color_data <= "111111100111";
      when "001001101000000" => color_data <= "111111100111";
      when "001001101000001" => color_data <= "111111100110";
      when "001001101000010" => color_data <= "111111010101";
      when "001001101000011" => color_data <= "111111100101";
      when "001001101000100" => color_data <= "111111100110";
      when "001001101000101" => color_data <= "111111100110";
      when "001001101000110" => color_data <= "111111101000";
      when "001001101000111" => color_data <= "111111111011";
      when "001001101001000" => color_data <= "111111101010";
      when "001001101001001" => color_data <= "111111101001";
      when "001001101001010" => color_data <= "111111111100";
      when "001001101001011" => color_data <= "111111100110";
      when "001001101001100" => color_data <= "111111000000";
      when "001001101001101" => color_data <= "111111010000";
      when "001001101001110" => color_data <= "111111010000";
      when "001001101001111" => color_data <= "111111010000";
      when "001001101010000" => color_data <= "100110000010";
      when "001001101010001" => color_data <= "001100110010";
      when "001001101010010" => color_data <= "100110000010";
      when "001001101010011" => color_data <= "110110100000";
      when "001001101010100" => color_data <= "111111000000";
      when "001001101010101" => color_data <= "110110100000";
      when "001001101010110" => color_data <= "101010000010";
      when "001001101010111" => color_data <= "000000000000";
      when "001001101011000" => color_data <= "000000000000";
      when "001001101011001" => color_data <= "000000000000";
      when "001001101011010" => color_data <= "000000000000";
      when "001001101011011" => color_data <= "001000100001";
      when "001001101011100" => color_data <= "111110110000";
      when "001001101011101" => color_data <= "111111000000";
      when "001001101011110" => color_data <= "110110100000";
      when "001001101011111" => color_data <= "000100010001";
      when "001001101100000" => color_data <= "000000000000";
      when "001001101100001" => color_data <= "000000000000";
      when "001001101100010" => color_data <= "000000000000";
      when "001001101100011" => color_data <= "000000000000";
      when "001001110000000" => color_data <= "000000000000";
      when "001001110000001" => color_data <= "000000000000";
      when "001001110000010" => color_data <= "000000000000";
      when "001001110000011" => color_data <= "000000000000";
      when "001001110000100" => color_data <= "000000000000";
      when "001001110000101" => color_data <= "000000000000";
      when "001001110000110" => color_data <= "000000000000";
      when "001001110000111" => color_data <= "000000000000";
      when "001001110001000" => color_data <= "011001010011";
      when "001001110001001" => color_data <= "111110110000";
      when "001001110001010" => color_data <= "111111000000";
      when "001001110001011" => color_data <= "100110000010";
      when "001001110001100" => color_data <= "000000000000";
      when "001001110001101" => color_data <= "000000000000";
      when "001001110001110" => color_data <= "000000000000";
      when "001001110001111" => color_data <= "000000000000";
      when "001001110010000" => color_data <= "000000000000";
      when "001001110010001" => color_data <= "001100110010";
      when "001001110010010" => color_data <= "110110010000";
      when "001001110010011" => color_data <= "111111000000";
      when "001001110010100" => color_data <= "111111010001";
      when "001001110010101" => color_data <= "111111010001";
      when "001001110010110" => color_data <= "111111010000";
      when "001001110010111" => color_data <= "111111010001";
      when "001001110011000" => color_data <= "111111111010";
      when "001001110011001" => color_data <= "111111111011";
      when "001001110011010" => color_data <= "111111101001";
      when "001001110011011" => color_data <= "111111101010";
      when "001001110011100" => color_data <= "111111101010";
      when "001001110011101" => color_data <= "111111101010";
      when "001001110011110" => color_data <= "111111101010";
      when "001001110011111" => color_data <= "111111101010";
      when "001001110100000" => color_data <= "111111101010";
      when "001001110100001" => color_data <= "111111101010";
      when "001001110100010" => color_data <= "111111101010";
      when "001001110100011" => color_data <= "111111111010";
      when "001001110100100" => color_data <= "111111101010";
      when "001001110100101" => color_data <= "111111101001";
      when "001001110100110" => color_data <= "111111101001";
      when "001001110100111" => color_data <= "111111100101";
      when "001001110101000" => color_data <= "111111000000";
      when "001001110101001" => color_data <= "111111010000";
      when "001001110101010" => color_data <= "111111010001";
      when "001001110101011" => color_data <= "111111010000";
      when "001001110101100" => color_data <= "111111010000";
      when "001001110101101" => color_data <= "111111010000";
      when "001001110101110" => color_data <= "111111010000";
      when "001001110101111" => color_data <= "111111010000";
      when "001001110110000" => color_data <= "111111010000";
      when "001001110110001" => color_data <= "111111010000";
      when "001001110110010" => color_data <= "111111010000";
      when "001001110110011" => color_data <= "111111010000";
      when "001001110110100" => color_data <= "111111010000";
      when "001001110110101" => color_data <= "111111010000";
      when "001001110110110" => color_data <= "111111010000";
      when "001001110110111" => color_data <= "111111010000";
      when "001001110111000" => color_data <= "111111010000";
      when "001001110111001" => color_data <= "111111010000";
      when "001001110111010" => color_data <= "111111010000";
      when "001001110111011" => color_data <= "111111010000";
      when "001001110111100" => color_data <= "111111010000";
      when "001001110111101" => color_data <= "111111010000";
      when "001001110111110" => color_data <= "111111010011";
      when "001001110111111" => color_data <= "111111100110";
      when "001001111000000" => color_data <= "111111010101";
      when "001001111000001" => color_data <= "111111100101";
      when "001001111000010" => color_data <= "111111100110";
      when "001001111000011" => color_data <= "111111101000";
      when "001001111000100" => color_data <= "111111101010";
      when "001001111000101" => color_data <= "111111111011";
      when "001001111000110" => color_data <= "111111101010";
      when "001001111000111" => color_data <= "111111101001";
      when "001001111001000" => color_data <= "111111101001";
      when "001001111001001" => color_data <= "111111101010";
      when "001001111001010" => color_data <= "111111111010";
      when "001001111001011" => color_data <= "111111111011";
      when "001001111001100" => color_data <= "111111010010";
      when "001001111001101" => color_data <= "111111010000";
      when "001001111001110" => color_data <= "111111010000";
      when "001001111001111" => color_data <= "111111010000";
      when "001001111010000" => color_data <= "111111000000";
      when "001001111010001" => color_data <= "111110110000";
      when "001001111010010" => color_data <= "111110110000";
      when "001001111010011" => color_data <= "111111000001";
      when "001001111010100" => color_data <= "111110110000";
      when "001001111010101" => color_data <= "110110100000";
      when "001001111010110" => color_data <= "000000000000";
      when "001001111010111" => color_data <= "000000000000";
      when "001001111011000" => color_data <= "000000000000";
      when "001001111011001" => color_data <= "000000000000";
      when "001001111011010" => color_data <= "000000000000";
      when "001001111011011" => color_data <= "010101000010";
      when "001001111011100" => color_data <= "111110110000";
      when "001001111011101" => color_data <= "111111000000";
      when "001001111011110" => color_data <= "101010000010";
      when "001001111011111" => color_data <= "000000000000";
      when "001001111100000" => color_data <= "000000000000";
      when "001001111100001" => color_data <= "000000000000";
      when "001001111100010" => color_data <= "000000000000";
      when "001001111100011" => color_data <= "000000000000";
      when "001010000000000" => color_data <= "000000000000";
      when "001010000000001" => color_data <= "000000000000";
      when "001010000000010" => color_data <= "000000000000";
      when "001010000000011" => color_data <= "000000000000";
      when "001010000000100" => color_data <= "000000000000";
      when "001010000000101" => color_data <= "000000000000";
      when "001010000000110" => color_data <= "000000000000";
      when "001010000000111" => color_data <= "000000000000";
      when "001010000001000" => color_data <= "001100110010";
      when "001010000001001" => color_data <= "110110100000";
      when "001010000001010" => color_data <= "111111000000";
      when "001010000001011" => color_data <= "110010010001";
      when "001010000001100" => color_data <= "000000000000";
      when "001010000001101" => color_data <= "000000000000";
      when "001010000001110" => color_data <= "000000000000";
      when "001010000001111" => color_data <= "000000000000";
      when "001010000010000" => color_data <= "000000000000";
      when "001010000010001" => color_data <= "000000000000";
      when "001010000010010" => color_data <= "010001000010";
      when "001010000010011" => color_data <= "110110100000";
      when "001010000010100" => color_data <= "111111010000";
      when "001010000010101" => color_data <= "111111010000";
      when "001010000010110" => color_data <= "111111010000";
      when "001010000010111" => color_data <= "111111101000";
      when "001010000011000" => color_data <= "111111111011";
      when "001010000011001" => color_data <= "111111101001";
      when "001010000011010" => color_data <= "111111101010";
      when "001010000011011" => color_data <= "111111101010";
      when "001010000011100" => color_data <= "111111101010";
      when "001010000011101" => color_data <= "111111101010";
      when "001010000011110" => color_data <= "111111101010";
      when "001010000011111" => color_data <= "111111101010";
      when "001010000100000" => color_data <= "111111101010";
      when "001010000100001" => color_data <= "111111101010";
      when "001010000100010" => color_data <= "111111101010";
      when "001010000100011" => color_data <= "111111101010";
      when "001010000100100" => color_data <= "111111101010";
      when "001010000100101" => color_data <= "111111101010";
      when "001010000100110" => color_data <= "111111111010";
      when "001010000100111" => color_data <= "111111101001";
      when "001010000101000" => color_data <= "111111010001";
      when "001010000101001" => color_data <= "111111010000";
      when "001010000101010" => color_data <= "111111010000";
      when "001010000101011" => color_data <= "111111010000";
      when "001010000101100" => color_data <= "111111010000";
      when "001010000101101" => color_data <= "111111010000";
      when "001010000101110" => color_data <= "111111010000";
      when "001010000101111" => color_data <= "111111010000";
      when "001010000110000" => color_data <= "111111010000";
      when "001010000110001" => color_data <= "111111010000";
      when "001010000110010" => color_data <= "111111010000";
      when "001010000110011" => color_data <= "111111010000";
      when "001010000110100" => color_data <= "111111010000";
      when "001010000110101" => color_data <= "111111010000";
      when "001010000110110" => color_data <= "111111010000";
      when "001010000110111" => color_data <= "111111010000";
      when "001010000111000" => color_data <= "111111010000";
      when "001010000111001" => color_data <= "111111010000";
      when "001010000111010" => color_data <= "111111010000";
      when "001010000111011" => color_data <= "111111010000";
      when "001010000111100" => color_data <= "111111010000";
      when "001010000111101" => color_data <= "111111010000";
      when "001010000111110" => color_data <= "111111010000";
      when "001010000111111" => color_data <= "111111100100";
      when "001010001000000" => color_data <= "111111101000";
      when "001010001000001" => color_data <= "111111101001";
      when "001010001000010" => color_data <= "111111111010";
      when "001010001000011" => color_data <= "111111111010";
      when "001010001000100" => color_data <= "111111101010";
      when "001010001000101" => color_data <= "111111101001";
      when "001010001000110" => color_data <= "111111101010";
      when "001010001000111" => color_data <= "111111101010";
      when "001010001001000" => color_data <= "111111101001";
      when "001010001001001" => color_data <= "111111101010";
      when "001010001001010" => color_data <= "111111101001";
      when "001010001001011" => color_data <= "111111111011";
      when "001010001001100" => color_data <= "111111101000";
      when "001010001001101" => color_data <= "111111010000";
      when "001010001001110" => color_data <= "111111010000";
      when "001010001001111" => color_data <= "111111010000";
      when "001010001010000" => color_data <= "111111010000";
      when "001010001010001" => color_data <= "111111000001";
      when "001010001010010" => color_data <= "111111000001";
      when "001010001010011" => color_data <= "111110110000";
      when "001010001010100" => color_data <= "110110100000";
      when "001010001010101" => color_data <= "001000100001";
      when "001010001010110" => color_data <= "000000000000";
      when "001010001010111" => color_data <= "000000000000";
      when "001010001011000" => color_data <= "000000000000";
      when "001010001011001" => color_data <= "000000000000";
      when "001010001011010" => color_data <= "000000000000";
      when "001010001011011" => color_data <= "100001110010";
      when "001010001011100" => color_data <= "111110110000";
      when "001010001011101" => color_data <= "111110110000";
      when "001010001011110" => color_data <= "100001110010";
      when "001010001011111" => color_data <= "000000000000";
      when "001010001100000" => color_data <= "000000000000";
      when "001010001100001" => color_data <= "000000000000";
      when "001010001100010" => color_data <= "000000000000";
      when "001010001100011" => color_data <= "000000000000";
      when "001010010000000" => color_data <= "000000000000";
      when "001010010000001" => color_data <= "000000000000";
      when "001010010000010" => color_data <= "000000000000";
      when "001010010000011" => color_data <= "000000000000";
      when "001010010000100" => color_data <= "000000000000";
      when "001010010000101" => color_data <= "000000000000";
      when "001010010000110" => color_data <= "000000000000";
      when "001010010000111" => color_data <= "000000000000";
      when "001010010001000" => color_data <= "000000000000";
      when "001010010001001" => color_data <= "110010010000";
      when "001010010001010" => color_data <= "111111000000";
      when "001010010001011" => color_data <= "110110100000";
      when "001010010001100" => color_data <= "010001000010";
      when "001010010001101" => color_data <= "000000000000";
      when "001010010001110" => color_data <= "000000000000";
      when "001010010001111" => color_data <= "000000000000";
      when "001010010010000" => color_data <= "000000000000";
      when "001010010010001" => color_data <= "000000000000";
      when "001010010010010" => color_data <= "000000000000";
      when "001010010010011" => color_data <= "001000100001";
      when "001010010010100" => color_data <= "110110110000";
      when "001010010010101" => color_data <= "111111000000";
      when "001010010010110" => color_data <= "111111100110";
      when "001010010010111" => color_data <= "111111111100";
      when "001010010011000" => color_data <= "111111101001";
      when "001010010011001" => color_data <= "111111101010";
      when "001010010011010" => color_data <= "111111101010";
      when "001010010011011" => color_data <= "111111101010";
      when "001010010011100" => color_data <= "111111101010";
      when "001010010011101" => color_data <= "111111101010";
      when "001010010011110" => color_data <= "111111101010";
      when "001010010011111" => color_data <= "111111101010";
      when "001010010100000" => color_data <= "111111101010";
      when "001010010100001" => color_data <= "111111101010";
      when "001010010100010" => color_data <= "111111101010";
      when "001010010100011" => color_data <= "111111101010";
      when "001010010100100" => color_data <= "111111101010";
      when "001010010100101" => color_data <= "111111101001";
      when "001010010100110" => color_data <= "111111101010";
      when "001010010100111" => color_data <= "111111111011";
      when "001010010101000" => color_data <= "111111010011";
      when "001010010101001" => color_data <= "111111010000";
      when "001010010101010" => color_data <= "111111010000";
      when "001010010101011" => color_data <= "111111010000";
      when "001010010101100" => color_data <= "111111010000";
      when "001010010101101" => color_data <= "111111010000";
      when "001010010101110" => color_data <= "111111010000";
      when "001010010101111" => color_data <= "111111010000";
      when "001010010110000" => color_data <= "111111010000";
      when "001010010110001" => color_data <= "111111010001";
      when "001010010110010" => color_data <= "111111010000";
      when "001010010110011" => color_data <= "111111010000";
      when "001010010110100" => color_data <= "111111010000";
      when "001010010110101" => color_data <= "111111010001";
      when "001010010110110" => color_data <= "111111010000";
      when "001010010110111" => color_data <= "111111010000";
      when "001010010111000" => color_data <= "111111010000";
      when "001010010111001" => color_data <= "111111010000";
      when "001010010111010" => color_data <= "111111010000";
      when "001010010111011" => color_data <= "111111010000";
      when "001010010111100" => color_data <= "111111010000";
      when "001010010111101" => color_data <= "111111010000";
      when "001010010111110" => color_data <= "111111010000";
      when "001010010111111" => color_data <= "111111101001";
      when "001010011000000" => color_data <= "111111111011";
      when "001010011000001" => color_data <= "111111101010";
      when "001010011000010" => color_data <= "111111101010";
      when "001010011000011" => color_data <= "111111101001";
      when "001010011000100" => color_data <= "111111101010";
      when "001010011000101" => color_data <= "111111101010";
      when "001010011000110" => color_data <= "111111101010";
      when "001010011000111" => color_data <= "111111101010";
      when "001010011001000" => color_data <= "111111101010";
      when "001010011001001" => color_data <= "111111101010";
      when "001010011001010" => color_data <= "111111101010";
      when "001010011001011" => color_data <= "111111101010";
      when "001010011001100" => color_data <= "111111111011";
      when "001010011001101" => color_data <= "111111010100";
      when "001010011001110" => color_data <= "111111000000";
      when "001010011001111" => color_data <= "111111010000";
      when "001010011010000" => color_data <= "111111010000";
      when "001010011010001" => color_data <= "111111000000";
      when "001010011010010" => color_data <= "111110110000";
      when "001010011010011" => color_data <= "110010100000";
      when "001010011010100" => color_data <= "000100010001";
      when "001010011010101" => color_data <= "000000000000";
      when "001010011010110" => color_data <= "000000000000";
      when "001010011010111" => color_data <= "000000000000";
      when "001010011011000" => color_data <= "000000000000";
      when "001010011011001" => color_data <= "000000000000";
      when "001010011011010" => color_data <= "000000000000";
      when "001010011011011" => color_data <= "101110010001";
      when "001010011011100" => color_data <= "111111000000";
      when "001010011011101" => color_data <= "111110110000";
      when "001010011011110" => color_data <= "010101000010";
      when "001010011011111" => color_data <= "000000000000";
      when "001010011100000" => color_data <= "000000000000";
      when "001010011100001" => color_data <= "000000000000";
      when "001010011100010" => color_data <= "000000000000";
      when "001010011100011" => color_data <= "000000000000";
      when "001010100000000" => color_data <= "000000000000";
      when "001010100000001" => color_data <= "000000000000";
      when "001010100000010" => color_data <= "000000000000";
      when "001010100000011" => color_data <= "000000000000";
      when "001010100000100" => color_data <= "000000000000";
      when "001010100000101" => color_data <= "000000000000";
      when "001010100000110" => color_data <= "000000000000";
      when "001010100000111" => color_data <= "000000000000";
      when "001010100001000" => color_data <= "000000000000";
      when "001010100001001" => color_data <= "100001110010";
      when "001010100001010" => color_data <= "111110110000";
      when "001010100001011" => color_data <= "111110110000";
      when "001010100001100" => color_data <= "100001110010";
      when "001010100001101" => color_data <= "000000000000";
      when "001010100001110" => color_data <= "000000000000";
      when "001010100001111" => color_data <= "000000000000";
      when "001010100010000" => color_data <= "000000000000";
      when "001010100010001" => color_data <= "000000000000";
      when "001010100010010" => color_data <= "000000000000";
      when "001010100010011" => color_data <= "000000000000";
      when "001010100010100" => color_data <= "101010010010";
      when "001010100010101" => color_data <= "111111010010";
      when "001010100010110" => color_data <= "111111111010";
      when "001010100010111" => color_data <= "111111101010";
      when "001010100011000" => color_data <= "111111101001";
      when "001010100011001" => color_data <= "111111101010";
      when "001010100011010" => color_data <= "111111101010";
      when "001010100011011" => color_data <= "111111101010";
      when "001010100011100" => color_data <= "111111101010";
      when "001010100011101" => color_data <= "111111101010";
      when "001010100011110" => color_data <= "111111101010";
      when "001010100011111" => color_data <= "111111101010";
      when "001010100100000" => color_data <= "111111101010";
      when "001010100100001" => color_data <= "111111101010";
      when "001010100100010" => color_data <= "111111101010";
      when "001010100100011" => color_data <= "111111101010";
      when "001010100100100" => color_data <= "111111101010";
      when "001010100100101" => color_data <= "111111101010";
      when "001010100100110" => color_data <= "111111101010";
      when "001010100100111" => color_data <= "111111111011";
      when "001010100101000" => color_data <= "111111100101";
      when "001010100101001" => color_data <= "111111000000";
      when "001010100101010" => color_data <= "111111010000";
      when "001010100101011" => color_data <= "111111010000";
      when "001010100101100" => color_data <= "111111010000";
      when "001010100101101" => color_data <= "111111010000";
      when "001010100101110" => color_data <= "111111010000";
      when "001010100101111" => color_data <= "111111010000";
      when "001010100110000" => color_data <= "111111010000";
      when "001010100110001" => color_data <= "111111010000";
      when "001010100110010" => color_data <= "111111010010";
      when "001010100110011" => color_data <= "111111100101";
      when "001010100110100" => color_data <= "111111010001";
      when "001010100110101" => color_data <= "111111010000";
      when "001010100110110" => color_data <= "111111010000";
      when "001010100110111" => color_data <= "111111010000";
      when "001010100111000" => color_data <= "111111010000";
      when "001010100111001" => color_data <= "111111010000";
      when "001010100111010" => color_data <= "111111010000";
      when "001010100111011" => color_data <= "111111010000";
      when "001010100111100" => color_data <= "111111010000";
      when "001010100111101" => color_data <= "111111000000";
      when "001010100111110" => color_data <= "111111010011";
      when "001010100111111" => color_data <= "111111111011";
      when "001010101000000" => color_data <= "111111101010";
      when "001010101000001" => color_data <= "111111101010";
      when "001010101000010" => color_data <= "111111101010";
      when "001010101000011" => color_data <= "111111101010";
      when "001010101000100" => color_data <= "111111101010";
      when "001010101000101" => color_data <= "111111101010";
      when "001010101000110" => color_data <= "111111101010";
      when "001010101000111" => color_data <= "111111101010";
      when "001010101001000" => color_data <= "111111101010";
      when "001010101001001" => color_data <= "111111101010";
      when "001010101001010" => color_data <= "111111101010";
      when "001010101001011" => color_data <= "111111101001";
      when "001010101001100" => color_data <= "111111111011";
      when "001010101001101" => color_data <= "111111101001";
      when "001010101001110" => color_data <= "111111010000";
      when "001010101001111" => color_data <= "111111010000";
      when "001010101010000" => color_data <= "111111000000";
      when "001010101010001" => color_data <= "110110100000";
      when "001010101010010" => color_data <= "100101110010";
      when "001010101010011" => color_data <= "000000000000";
      when "001010101010100" => color_data <= "000000000000";
      when "001010101010101" => color_data <= "000000000000";
      when "001010101010110" => color_data <= "000000000000";
      when "001010101010111" => color_data <= "000000000000";
      when "001010101011000" => color_data <= "000000000000";
      when "001010101011001" => color_data <= "000000000000";
      when "001010101011010" => color_data <= "001100110010";
      when "001010101011011" => color_data <= "110110100000";
      when "001010101011100" => color_data <= "111111000000";
      when "001010101011101" => color_data <= "110010100000";
      when "001010101011110" => color_data <= "000000000000";
      when "001010101011111" => color_data <= "000000000000";
      when "001010101100000" => color_data <= "000000000000";
      when "001010101100001" => color_data <= "000000000000";
      when "001010101100010" => color_data <= "000000000000";
      when "001010101100011" => color_data <= "000000000000";
      when "001010110000000" => color_data <= "000000000000";
      when "001010110000001" => color_data <= "000000000000";
      when "001010110000010" => color_data <= "000000000000";
      when "001010110000011" => color_data <= "000000000000";
      when "001010110000100" => color_data <= "000000000000";
      when "001010110000101" => color_data <= "000000000000";
      when "001010110000110" => color_data <= "000000000000";
      when "001010110000111" => color_data <= "000000000000";
      when "001010110001000" => color_data <= "000000000000";
      when "001010110001001" => color_data <= "010001000010";
      when "001010110001010" => color_data <= "111110110000";
      when "001010110001011" => color_data <= "111111000000";
      when "001010110001100" => color_data <= "101110010001";
      when "001010110001101" => color_data <= "000000000000";
      when "001010110001110" => color_data <= "000000000000";
      when "001010110001111" => color_data <= "000000000000";
      when "001010110010000" => color_data <= "000000000000";
      when "001010110010001" => color_data <= "000000000000";
      when "001010110010010" => color_data <= "000000000000";
      when "001010110010011" => color_data <= "000000000000";
      when "001010110010100" => color_data <= "011001100011";
      when "001010110010101" => color_data <= "111111100101";
      when "001010110010110" => color_data <= "111111101010";
      when "001010110010111" => color_data <= "111111101010";
      when "001010110011000" => color_data <= "111111101010";
      when "001010110011001" => color_data <= "111111101010";
      when "001010110011010" => color_data <= "111111101010";
      when "001010110011011" => color_data <= "111111101010";
      when "001010110011100" => color_data <= "111111101010";
      when "001010110011101" => color_data <= "111111101010";
      when "001010110011110" => color_data <= "111111101010";
      when "001010110011111" => color_data <= "111111101010";
      when "001010110100000" => color_data <= "111111101010";
      when "001010110100001" => color_data <= "111111101010";
      when "001010110100010" => color_data <= "111111101010";
      when "001010110100011" => color_data <= "111111101010";
      when "001010110100100" => color_data <= "111111101010";
      when "001010110100101" => color_data <= "111111101010";
      when "001010110100110" => color_data <= "111111101010";
      when "001010110100111" => color_data <= "111111111011";
      when "001010110101000" => color_data <= "111111100111";
      when "001010110101001" => color_data <= "111111000000";
      when "001010110101010" => color_data <= "111111010000";
      when "001010110101011" => color_data <= "111111010000";
      when "001010110101100" => color_data <= "111111010000";
      when "001010110101101" => color_data <= "111111010000";
      when "001010110101110" => color_data <= "111111010000";
      when "001010110101111" => color_data <= "111111010000";
      when "001010110110000" => color_data <= "111111010000";
      when "001010110110001" => color_data <= "111111010000";
      when "001010110110010" => color_data <= "111111010010";
      when "001010110110011" => color_data <= "111111101001";
      when "001010110110100" => color_data <= "111111010100";
      when "001010110110101" => color_data <= "111111010000";
      when "001010110110110" => color_data <= "111111010000";
      when "001010110110111" => color_data <= "111111010000";
      when "001010110111000" => color_data <= "111111010000";
      when "001010110111001" => color_data <= "111111010000";
      when "001010110111010" => color_data <= "111111010000";
      when "001010110111011" => color_data <= "111111010000";
      when "001010110111100" => color_data <= "111111010000";
      when "001010110111101" => color_data <= "111111000000";
      when "001010110111110" => color_data <= "111111100110";
      when "001010110111111" => color_data <= "111111111011";
      when "001010111000000" => color_data <= "111111101010";
      when "001010111000001" => color_data <= "111111101001";
      when "001010111000010" => color_data <= "111111101010";
      when "001010111000011" => color_data <= "111111101010";
      when "001010111000100" => color_data <= "111111101010";
      when "001010111000101" => color_data <= "111111101010";
      when "001010111000110" => color_data <= "111111101010";
      when "001010111000111" => color_data <= "111111101010";
      when "001010111001000" => color_data <= "111111101010";
      when "001010111001001" => color_data <= "111111101010";
      when "001010111001010" => color_data <= "111111101010";
      when "001010111001011" => color_data <= "111111101010";
      when "001010111001100" => color_data <= "111111101001";
      when "001010111001101" => color_data <= "111111111011";
      when "001010111001110" => color_data <= "111111100101";
      when "001010111001111" => color_data <= "111111010000";
      when "001010111010000" => color_data <= "100101110010";
      when "001010111010001" => color_data <= "001100110010";
      when "001010111010010" => color_data <= "000000000000";
      when "001010111010011" => color_data <= "000000000000";
      when "001010111010100" => color_data <= "000000000000";
      when "001010111010101" => color_data <= "000000000000";
      when "001010111010110" => color_data <= "000000000000";
      when "001010111010111" => color_data <= "000000000000";
      when "001010111011000" => color_data <= "000000000000";
      when "001010111011001" => color_data <= "000000000000";
      when "001010111011010" => color_data <= "011101100011";
      when "001010111011011" => color_data <= "111110110000";
      when "001010111011100" => color_data <= "111110110000";
      when "001010111011101" => color_data <= "100110000010";
      when "001010111011110" => color_data <= "000000000000";
      when "001010111011111" => color_data <= "000000000000";
      when "001010111100000" => color_data <= "000000000000";
      when "001010111100001" => color_data <= "000000000000";
      when "001010111100010" => color_data <= "000000000000";
      when "001010111100011" => color_data <= "000000000000";
      when "001011000000000" => color_data <= "000000000000";
      when "001011000000001" => color_data <= "000000000000";
      when "001011000000010" => color_data <= "000000000000";
      when "001011000000011" => color_data <= "000000000000";
      when "001011000000100" => color_data <= "000000000000";
      when "001011000000101" => color_data <= "000000000000";
      when "001011000000110" => color_data <= "000000000000";
      when "001011000000111" => color_data <= "000000000000";
      when "001011000001000" => color_data <= "000000000000";
      when "001011000001001" => color_data <= "000000000000";
      when "001011000001010" => color_data <= "110110100000";
      when "001011000001011" => color_data <= "111111000000";
      when "001011000001100" => color_data <= "101110010001";
      when "001011000001101" => color_data <= "000000000000";
      when "001011000001110" => color_data <= "000000000000";
      when "001011000001111" => color_data <= "000000000000";
      when "001011000010000" => color_data <= "000000000000";
      when "001011000010001" => color_data <= "000000000000";
      when "001011000010010" => color_data <= "000000000000";
      when "001011000010011" => color_data <= "000000000000";
      when "001011000010100" => color_data <= "010001000010";
      when "001011000010101" => color_data <= "111111010100";
      when "001011000010110" => color_data <= "111111101001";
      when "001011000010111" => color_data <= "111111101010";
      when "001011000011000" => color_data <= "111111101010";
      when "001011000011001" => color_data <= "111111101010";
      when "001011000011010" => color_data <= "111111101010";
      when "001011000011011" => color_data <= "111111101010";
      when "001011000011100" => color_data <= "111111101010";
      when "001011000011101" => color_data <= "111111101010";
      when "001011000011110" => color_data <= "111111101010";
      when "001011000011111" => color_data <= "111111101010";
      when "001011000100000" => color_data <= "111111101010";
      when "001011000100001" => color_data <= "111111101010";
      when "001011000100010" => color_data <= "111111101010";
      when "001011000100011" => color_data <= "111111101010";
      when "001011000100100" => color_data <= "111111101010";
      when "001011000100101" => color_data <= "111111101010";
      when "001011000100110" => color_data <= "111111101010";
      when "001011000100111" => color_data <= "111111111010";
      when "001011000101000" => color_data <= "111111101001";
      when "001011000101001" => color_data <= "111111010001";
      when "001011000101010" => color_data <= "111111010000";
      when "001011000101011" => color_data <= "111111010000";
      when "001011000101100" => color_data <= "111111010000";
      when "001011000101101" => color_data <= "111111010000";
      when "001011000101110" => color_data <= "111111010000";
      when "001011000101111" => color_data <= "111111010000";
      when "001011000110000" => color_data <= "111111010000";
      when "001011000110001" => color_data <= "111111010000";
      when "001011000110010" => color_data <= "111111010011";
      when "001011000110011" => color_data <= "111111101010";
      when "001011000110100" => color_data <= "111111010100";
      when "001011000110101" => color_data <= "111111010000";
      when "001011000110110" => color_data <= "111111010000";
      when "001011000110111" => color_data <= "111111010000";
      when "001011000111000" => color_data <= "111111010000";
      when "001011000111001" => color_data <= "111111010000";
      when "001011000111010" => color_data <= "111111010000";
      when "001011000111011" => color_data <= "111111010000";
      when "001011000111100" => color_data <= "111111010000";
      when "001011000111101" => color_data <= "111111010001";
      when "001011000111110" => color_data <= "111111101010";
      when "001011000111111" => color_data <= "111111101010";
      when "001011001000000" => color_data <= "111111101010";
      when "001011001000001" => color_data <= "111111101010";
      when "001011001000010" => color_data <= "111111101010";
      when "001011001000011" => color_data <= "111111101010";
      when "001011001000100" => color_data <= "111111101010";
      when "001011001000101" => color_data <= "111111101010";
      when "001011001000110" => color_data <= "111111101010";
      when "001011001000111" => color_data <= "111111101010";
      when "001011001001000" => color_data <= "111111101010";
      when "001011001001001" => color_data <= "111111101010";
      when "001011001001010" => color_data <= "111111101010";
      when "001011001001011" => color_data <= "111111101010";
      when "001011001001100" => color_data <= "111111101001";
      when "001011001001101" => color_data <= "111111111011";
      when "001011001001110" => color_data <= "111111100111";
      when "001011001001111" => color_data <= "111111010010";
      when "001011001010000" => color_data <= "001000100001";
      when "001011001010001" => color_data <= "000000000000";
      when "001011001010010" => color_data <= "000000000000";
      when "001011001010011" => color_data <= "000000000000";
      when "001011001010100" => color_data <= "000000000000";
      when "001011001010101" => color_data <= "000000000000";
      when "001011001010110" => color_data <= "000000000000";
      when "001011001010111" => color_data <= "000000000000";
      when "001011001011000" => color_data <= "000000000000";
      when "001011001011001" => color_data <= "000000000000";
      when "001011001011010" => color_data <= "101010000010";
      when "001011001011011" => color_data <= "111111000000";
      when "001011001011100" => color_data <= "111110110000";
      when "001011001011101" => color_data <= "010101010011";
      when "001011001011110" => color_data <= "000000000000";
      when "001011001011111" => color_data <= "000000000000";
      when "001011001100000" => color_data <= "000000000000";
      when "001011001100001" => color_data <= "000000000000";
      when "001011001100010" => color_data <= "000000000000";
      when "001011001100011" => color_data <= "000000000000";
      when "001011010000000" => color_data <= "000000000000";
      when "001011010000001" => color_data <= "000000000000";
      when "001011010000010" => color_data <= "000000000000";
      when "001011010000011" => color_data <= "000000000000";
      when "001011010000100" => color_data <= "000000000000";
      when "001011010000101" => color_data <= "000000000000";
      when "001011010000110" => color_data <= "000000000000";
      when "001011010000111" => color_data <= "000000000000";
      when "001011010001000" => color_data <= "000000000000";
      when "001011010001001" => color_data <= "000000000000";
      when "001011010001010" => color_data <= "100001110010";
      when "001011010001011" => color_data <= "111110110000";
      when "001011010001100" => color_data <= "111111000001";
      when "001011010001101" => color_data <= "011001010011";
      when "001011010001110" => color_data <= "000000000000";
      when "001011010001111" => color_data <= "000000000000";
      when "001011010010000" => color_data <= "000000000000";
      when "001011010010001" => color_data <= "000000000000";
      when "001011010010010" => color_data <= "000000000000";
      when "001011010010011" => color_data <= "000000000000";
      when "001011010010100" => color_data <= "001100100010";
      when "001011010010101" => color_data <= "111111010011";
      when "001011010010110" => color_data <= "111111101000";
      when "001011010010111" => color_data <= "111111111010";
      when "001011010011000" => color_data <= "111111101010";
      when "001011010011001" => color_data <= "111111101010";
      when "001011010011010" => color_data <= "111111101010";
      when "001011010011011" => color_data <= "111111101010";
      when "001011010011100" => color_data <= "111111101010";
      when "001011010011101" => color_data <= "111111101010";
      when "001011010011110" => color_data <= "111111101010";
      when "001011010011111" => color_data <= "111111101010";
      when "001011010100000" => color_data <= "111111101010";
      when "001011010100001" => color_data <= "111111101010";
      when "001011010100010" => color_data <= "111111101010";
      when "001011010100011" => color_data <= "111111101010";
      when "001011010100100" => color_data <= "111111101010";
      when "001011010100101" => color_data <= "111111101010";
      when "001011010100110" => color_data <= "111111101010";
      when "001011010100111" => color_data <= "111111101010";
      when "001011010101000" => color_data <= "111111111011";
      when "001011010101001" => color_data <= "111111010011";
      when "001011010101010" => color_data <= "111111010000";
      when "001011010101011" => color_data <= "111111010000";
      when "001011010101100" => color_data <= "111111010000";
      when "001011010101101" => color_data <= "111111010000";
      when "001011010101110" => color_data <= "111111010000";
      when "001011010101111" => color_data <= "111111010000";
      when "001011010110000" => color_data <= "111111010000";
      when "001011010110001" => color_data <= "111111010000";
      when "001011010110010" => color_data <= "111111010010";
      when "001011010110011" => color_data <= "111111100101";
      when "001011010110100" => color_data <= "111111010001";
      when "001011010110101" => color_data <= "111111010000";
      when "001011010110110" => color_data <= "111111010000";
      when "001011010110111" => color_data <= "111111010000";
      when "001011010111000" => color_data <= "111111010000";
      when "001011010111001" => color_data <= "111111010000";
      when "001011010111010" => color_data <= "111111010000";
      when "001011010111011" => color_data <= "111111010000";
      when "001011010111100" => color_data <= "111111010000";
      when "001011010111101" => color_data <= "111111010100";
      when "001011010111110" => color_data <= "111111111011";
      when "001011010111111" => color_data <= "111111101010";
      when "001011011000000" => color_data <= "111111101010";
      when "001011011000001" => color_data <= "111111101010";
      when "001011011000010" => color_data <= "111111101010";
      when "001011011000011" => color_data <= "111111101010";
      when "001011011000100" => color_data <= "111111101010";
      when "001011011000101" => color_data <= "111111101010";
      when "001011011000110" => color_data <= "111111101010";
      when "001011011000111" => color_data <= "111111101010";
      when "001011011001000" => color_data <= "111111101010";
      when "001011011001001" => color_data <= "111111101010";
      when "001011011001010" => color_data <= "111111101010";
      when "001011011001011" => color_data <= "111111101001";
      when "001011011001100" => color_data <= "111111101010";
      when "001011011001101" => color_data <= "111111101010";
      when "001011011001110" => color_data <= "111111100101";
      when "001011011001111" => color_data <= "100001110010";
      when "001011011010000" => color_data <= "000000000000";
      when "001011011010001" => color_data <= "000000000000";
      when "001011011010010" => color_data <= "000000000000";
      when "001011011010011" => color_data <= "000000000000";
      when "001011011010100" => color_data <= "000000000000";
      when "001011011010101" => color_data <= "000000000000";
      when "001011011010110" => color_data <= "000000000000";
      when "001011011010111" => color_data <= "000000000000";
      when "001011011011000" => color_data <= "000000000000";
      when "001011011011001" => color_data <= "001000100001";
      when "001011011011010" => color_data <= "110110100000";
      when "001011011011011" => color_data <= "111111000000";
      when "001011011011100" => color_data <= "110110100000";
      when "001011011011101" => color_data <= "000000000000";
      when "001011011011110" => color_data <= "000000000000";
      when "001011011011111" => color_data <= "000000000000";
      when "001011011100000" => color_data <= "000000000000";
      when "001011011100001" => color_data <= "000000000000";
      when "001011011100010" => color_data <= "000000000000";
      when "001011011100011" => color_data <= "000000000000";
      when "001011100000000" => color_data <= "000000000000";
      when "001011100000001" => color_data <= "000000000000";
      when "001011100000010" => color_data <= "000000000000";
      when "001011100000011" => color_data <= "000000000000";
      when "001011100000100" => color_data <= "000000000000";
      when "001011100000101" => color_data <= "000000000000";
      when "001011100000110" => color_data <= "000000000000";
      when "001011100000111" => color_data <= "000000000000";
      when "001011100001000" => color_data <= "000000000000";
      when "001011100001001" => color_data <= "000000000000";
      when "001011100001010" => color_data <= "001100110010";
      when "001011100001011" => color_data <= "110110100000";
      when "001011100001100" => color_data <= "111111000000";
      when "001011100001101" => color_data <= "110110100000";
      when "001011100001110" => color_data <= "000100010001";
      when "001011100001111" => color_data <= "000000000000";
      when "001011100010000" => color_data <= "000000000000";
      when "001011100010001" => color_data <= "000000000000";
      when "001011100010010" => color_data <= "000000000000";
      when "001011100010011" => color_data <= "000000000000";
      when "001011100010100" => color_data <= "000100010001";
      when "001011100010101" => color_data <= "101010010010";
      when "001011100010110" => color_data <= "111111100110";
      when "001011100010111" => color_data <= "111111111010";
      when "001011100011000" => color_data <= "111111101010";
      when "001011100011001" => color_data <= "111111101010";
      when "001011100011010" => color_data <= "111111101010";
      when "001011100011011" => color_data <= "111111101010";
      when "001011100011100" => color_data <= "111111101010";
      when "001011100011101" => color_data <= "111111101010";
      when "001011100011110" => color_data <= "111111101010";
      when "001011100011111" => color_data <= "111111101010";
      when "001011100100000" => color_data <= "111111101010";
      when "001011100100001" => color_data <= "111111101010";
      when "001011100100010" => color_data <= "111111101010";
      when "001011100100011" => color_data <= "111111101010";
      when "001011100100100" => color_data <= "111111101010";
      when "001011100100101" => color_data <= "111111101010";
      when "001011100100110" => color_data <= "111111101010";
      when "001011100100111" => color_data <= "111111101010";
      when "001011100101000" => color_data <= "111111111011";
      when "001011100101001" => color_data <= "111111100101";
      when "001011100101010" => color_data <= "111111010000";
      when "001011100101011" => color_data <= "111111010000";
      when "001011100101100" => color_data <= "111111010000";
      when "001011100101101" => color_data <= "111111010000";
      when "001011100101110" => color_data <= "111111010000";
      when "001011100101111" => color_data <= "111111010000";
      when "001011100110000" => color_data <= "111111010000";
      when "001011100110001" => color_data <= "111111010001";
      when "001011100110010" => color_data <= "111111010000";
      when "001011100110011" => color_data <= "111111010000";
      when "001011100110100" => color_data <= "111111010000";
      when "001011100110101" => color_data <= "111111010001";
      when "001011100110110" => color_data <= "111111010000";
      when "001011100110111" => color_data <= "111111010000";
      when "001011100111000" => color_data <= "111111010000";
      when "001011100111001" => color_data <= "111111010000";
      when "001011100111010" => color_data <= "111111010000";
      when "001011100111011" => color_data <= "111111010000";
      when "001011100111100" => color_data <= "111111010000";
      when "001011100111101" => color_data <= "111111100111";
      when "001011100111110" => color_data <= "111111111011";
      when "001011100111111" => color_data <= "111111101001";
      when "001011101000000" => color_data <= "111111101010";
      when "001011101000001" => color_data <= "111111101010";
      when "001011101000010" => color_data <= "111111101010";
      when "001011101000011" => color_data <= "111111101010";
      when "001011101000100" => color_data <= "111111101010";
      when "001011101000101" => color_data <= "111111101010";
      when "001011101000110" => color_data <= "111111101010";
      when "001011101000111" => color_data <= "111111101010";
      when "001011101001000" => color_data <= "111111101010";
      when "001011101001001" => color_data <= "111111101010";
      when "001011101001010" => color_data <= "111111101010";
      when "001011101001011" => color_data <= "111111101010";
      when "001011101001100" => color_data <= "111111111010";
      when "001011101001101" => color_data <= "111111101000";
      when "001011101001110" => color_data <= "111111010100";
      when "001011101001111" => color_data <= "011001100011";
      when "001011101010000" => color_data <= "000000000000";
      when "001011101010001" => color_data <= "000000000000";
      when "001011101010010" => color_data <= "000000000000";
      when "001011101010011" => color_data <= "000000000000";
      when "001011101010100" => color_data <= "000000000000";
      when "001011101010101" => color_data <= "000000000000";
      when "001011101010110" => color_data <= "000000000000";
      when "001011101010111" => color_data <= "000000000000";
      when "001011101011000" => color_data <= "000000000000";
      when "001011101011001" => color_data <= "100110000010";
      when "001011101011010" => color_data <= "111110110000";
      when "001011101011011" => color_data <= "111110110000";
      when "001011101011100" => color_data <= "100110000010";
      when "001011101011101" => color_data <= "000000000000";
      when "001011101011110" => color_data <= "000000000000";
      when "001011101011111" => color_data <= "000000000000";
      when "001011101100000" => color_data <= "000000000000";
      when "001011101100001" => color_data <= "000000000000";
      when "001011101100010" => color_data <= "000000000000";
      when "001011101100011" => color_data <= "000000000000";
      when "001011110000000" => color_data <= "000000000000";
      when "001011110000001" => color_data <= "000000000000";
      when "001011110000010" => color_data <= "000000000000";
      when "001011110000011" => color_data <= "000000000000";
      when "001011110000100" => color_data <= "000000000000";
      when "001011110000101" => color_data <= "000000000000";
      when "001011110000110" => color_data <= "000000000000";
      when "001011110000111" => color_data <= "000000000000";
      when "001011110001000" => color_data <= "000000000000";
      when "001011110001001" => color_data <= "000000000000";
      when "001011110001010" => color_data <= "000000000000";
      when "001011110001011" => color_data <= "101110010001";
      when "001011110001100" => color_data <= "111110110000";
      when "001011110001101" => color_data <= "111110110000";
      when "001011110001110" => color_data <= "011101100011";
      when "001011110001111" => color_data <= "000000000000";
      when "001011110010000" => color_data <= "000000000000";
      when "001011110010001" => color_data <= "000000000000";
      when "001011110010010" => color_data <= "000000000000";
      when "001011110010011" => color_data <= "000000000000";
      when "001011110010100" => color_data <= "000000000000";
      when "001011110010101" => color_data <= "011101110011";
      when "001011110010110" => color_data <= "111111100101";
      when "001011110010111" => color_data <= "111111101010";
      when "001011110011000" => color_data <= "111111101001";
      when "001011110011001" => color_data <= "111111101010";
      when "001011110011010" => color_data <= "111111101010";
      when "001011110011011" => color_data <= "111111101010";
      when "001011110011100" => color_data <= "111111101010";
      when "001011110011101" => color_data <= "111111101010";
      when "001011110011110" => color_data <= "111111101010";
      when "001011110011111" => color_data <= "111111101010";
      when "001011110100000" => color_data <= "111111101010";
      when "001011110100001" => color_data <= "111111101010";
      when "001011110100010" => color_data <= "111111101010";
      when "001011110100011" => color_data <= "111111101010";
      when "001011110100100" => color_data <= "111111101010";
      when "001011110100101" => color_data <= "111111101010";
      when "001011110100110" => color_data <= "111111101010";
      when "001011110100111" => color_data <= "111111101010";
      when "001011110101000" => color_data <= "111111111011";
      when "001011110101001" => color_data <= "111111100111";
      when "001011110101010" => color_data <= "111111010000";
      when "001011110101011" => color_data <= "111111010000";
      when "001011110101100" => color_data <= "111111010001";
      when "001011110101101" => color_data <= "111111010000";
      when "001011110101110" => color_data <= "111111010000";
      when "001011110101111" => color_data <= "111111010000";
      when "001011110110000" => color_data <= "111111010000";
      when "001011110110001" => color_data <= "111111010000";
      when "001011110110010" => color_data <= "111111010000";
      when "001011110110011" => color_data <= "111111010000";
      when "001011110110100" => color_data <= "111111010000";
      when "001011110110101" => color_data <= "111111010000";
      when "001011110110110" => color_data <= "111111010000";
      when "001011110110111" => color_data <= "111111010000";
      when "001011110111000" => color_data <= "111111010000";
      when "001011110111001" => color_data <= "111111010000";
      when "001011110111010" => color_data <= "111111010000";
      when "001011110111011" => color_data <= "111111010000";
      when "001011110111100" => color_data <= "111111010010";
      when "001011110111101" => color_data <= "111111111010";
      when "001011110111110" => color_data <= "111111101010";
      when "001011110111111" => color_data <= "111111101010";
      when "001011111000000" => color_data <= "111111101010";
      when "001011111000001" => color_data <= "111111101010";
      when "001011111000010" => color_data <= "111111101010";
      when "001011111000011" => color_data <= "111111101010";
      when "001011111000100" => color_data <= "111111101010";
      when "001011111000101" => color_data <= "111111101010";
      when "001011111000110" => color_data <= "111111101010";
      when "001011111000111" => color_data <= "111111101010";
      when "001011111001000" => color_data <= "111111101010";
      when "001011111001001" => color_data <= "111111101010";
      when "001011111001010" => color_data <= "111111101010";
      when "001011111001011" => color_data <= "111111101001";
      when "001011111001100" => color_data <= "111111111011";
      when "001011111001101" => color_data <= "111111100111";
      when "001011111001110" => color_data <= "111111010100";
      when "001011111001111" => color_data <= "010101010010";
      when "001011111010000" => color_data <= "000000000000";
      when "001011111010001" => color_data <= "000000000000";
      when "001011111010010" => color_data <= "000000000000";
      when "001011111010011" => color_data <= "000000000000";
      when "001011111010100" => color_data <= "000000000000";
      when "001011111010101" => color_data <= "000000000000";
      when "001011111010110" => color_data <= "000000000000";
      when "001011111010111" => color_data <= "000000000000";
      when "001011111011000" => color_data <= "000000000000";
      when "001011111011001" => color_data <= "110110100000";
      when "001011111011010" => color_data <= "111111000000";
      when "001011111011011" => color_data <= "110110100000";
      when "001011111011100" => color_data <= "010000110010";
      when "001011111011101" => color_data <= "000000000000";
      when "001011111011110" => color_data <= "000000000000";
      when "001011111011111" => color_data <= "000000000000";
      when "001011111100000" => color_data <= "000000000000";
      when "001011111100001" => color_data <= "000000000000";
      when "001011111100010" => color_data <= "000000000000";
      when "001011111100011" => color_data <= "000000000000";
      when "001100000000000" => color_data <= "000000000000";
      when "001100000000001" => color_data <= "000000000000";
      when "001100000000010" => color_data <= "000000000000";
      when "001100000000011" => color_data <= "000000000000";
      when "001100000000100" => color_data <= "000000000000";
      when "001100000000101" => color_data <= "000000000000";
      when "001100000000110" => color_data <= "000000000000";
      when "001100000000111" => color_data <= "000000000000";
      when "001100000001000" => color_data <= "000000000000";
      when "001100000001001" => color_data <= "000000000000";
      when "001100000001010" => color_data <= "000000000000";
      when "001100000001011" => color_data <= "010101010010";
      when "001100000001100" => color_data <= "110110100000";
      when "001100000001101" => color_data <= "111111000000";
      when "001100000001110" => color_data <= "110110100000";
      when "001100000001111" => color_data <= "000000000000";
      when "001100000010000" => color_data <= "000000000000";
      when "001100000010001" => color_data <= "000000000000";
      when "001100000010010" => color_data <= "000000000000";
      when "001100000010011" => color_data <= "000000000000";
      when "001100000010100" => color_data <= "000000000000";
      when "001100000010101" => color_data <= "010001000010";
      when "001100000010110" => color_data <= "111111010011";
      when "001100000010111" => color_data <= "111111101000";
      when "001100000011000" => color_data <= "111111111010";
      when "001100000011001" => color_data <= "111111101010";
      when "001100000011010" => color_data <= "111111101010";
      when "001100000011011" => color_data <= "111111101010";
      when "001100000011100" => color_data <= "111111101010";
      when "001100000011101" => color_data <= "111111101010";
      when "001100000011110" => color_data <= "111111101010";
      when "001100000011111" => color_data <= "111111101010";
      when "001100000100000" => color_data <= "111111101010";
      when "001100000100001" => color_data <= "111111101010";
      when "001100000100010" => color_data <= "111111101010";
      when "001100000100011" => color_data <= "111111101010";
      when "001100000100100" => color_data <= "111111101010";
      when "001100000100101" => color_data <= "111111101010";
      when "001100000100110" => color_data <= "111111101010";
      when "001100000100111" => color_data <= "111111101001";
      when "001100000101000" => color_data <= "111111111010";
      when "001100000101001" => color_data <= "111111101001";
      when "001100000101010" => color_data <= "111111010001";
      when "001100000101011" => color_data <= "111111010000";
      when "001100000101100" => color_data <= "111111010000";
      when "001100000101101" => color_data <= "111111010000";
      when "001100000101110" => color_data <= "111111010000";
      when "001100000101111" => color_data <= "111111010000";
      when "001100000110000" => color_data <= "111111010000";
      when "001100000110001" => color_data <= "111111010000";
      when "001100000110010" => color_data <= "111111010000";
      when "001100000110011" => color_data <= "111111010000";
      when "001100000110100" => color_data <= "111111010000";
      when "001100000110101" => color_data <= "111111010000";
      when "001100000110110" => color_data <= "111111010000";
      when "001100000110111" => color_data <= "111111010000";
      when "001100000111000" => color_data <= "111111010000";
      when "001100000111001" => color_data <= "111111010000";
      when "001100000111010" => color_data <= "111111010000";
      when "001100000111011" => color_data <= "111111010000";
      when "001100000111100" => color_data <= "111111100110";
      when "001100000111101" => color_data <= "111111111011";
      when "001100000111110" => color_data <= "111111101001";
      when "001100000111111" => color_data <= "111111101010";
      when "001100001000000" => color_data <= "111111101010";
      when "001100001000001" => color_data <= "111111101010";
      when "001100001000010" => color_data <= "111111101010";
      when "001100001000011" => color_data <= "111111101010";
      when "001100001000100" => color_data <= "111111101010";
      when "001100001000101" => color_data <= "111111101010";
      when "001100001000110" => color_data <= "111111101010";
      when "001100001000111" => color_data <= "111111101010";
      when "001100001001000" => color_data <= "111111101010";
      when "001100001001001" => color_data <= "111111101010";
      when "001100001001010" => color_data <= "111111101010";
      when "001100001001011" => color_data <= "111111101010";
      when "001100001001100" => color_data <= "111111101010";
      when "001100001001101" => color_data <= "111111100110";
      when "001100001001110" => color_data <= "111111010100";
      when "001100001001111" => color_data <= "001100110010";
      when "001100001010000" => color_data <= "000000000000";
      when "001100001010001" => color_data <= "000000000000";
      when "001100001010010" => color_data <= "000000000000";
      when "001100001010011" => color_data <= "000000000000";
      when "001100001010100" => color_data <= "000000000000";
      when "001100001010101" => color_data <= "000000000000";
      when "001100001010110" => color_data <= "000000000000";
      when "001100001010111" => color_data <= "000000000000";
      when "001100001011000" => color_data <= "011101100011";
      when "001100001011001" => color_data <= "111110110000";
      when "001100001011010" => color_data <= "111111000000";
      when "001100001011011" => color_data <= "101110010001";
      when "001100001011100" => color_data <= "000000000000";
      when "001100001011101" => color_data <= "000000000000";
      when "001100001011110" => color_data <= "000000000000";
      when "001100001011111" => color_data <= "000000000000";
      when "001100001100000" => color_data <= "000000000000";
      when "001100001100001" => color_data <= "000000000000";
      when "001100001100010" => color_data <= "000000000000";
      when "001100001100011" => color_data <= "000000000000";
      when "001100010000000" => color_data <= "000000000000";
      when "001100010000001" => color_data <= "000000000000";
      when "001100010000010" => color_data <= "000000000000";
      when "001100010000011" => color_data <= "000000000000";
      when "001100010000100" => color_data <= "000000000000";
      when "001100010000101" => color_data <= "000000000000";
      when "001100010000110" => color_data <= "000000000000";
      when "001100010000111" => color_data <= "000000000000";
      when "001100010001000" => color_data <= "000000000000";
      when "001100010001001" => color_data <= "000000000000";
      when "001100010001010" => color_data <= "000000000000";
      when "001100010001011" => color_data <= "000000000000";
      when "001100010001100" => color_data <= "110110100000";
      when "001100010001101" => color_data <= "111111000000";
      when "001100010001110" => color_data <= "111110110000";
      when "001100010001111" => color_data <= "011001010011";
      when "001100010010000" => color_data <= "000000000000";
      when "001100010010001" => color_data <= "000000000000";
      when "001100010010010" => color_data <= "000000000000";
      when "001100010010011" => color_data <= "000000000000";
      when "001100010010100" => color_data <= "000000000000";
      when "001100010010101" => color_data <= "000100010001";
      when "001100010010110" => color_data <= "101110010001";
      when "001100010010111" => color_data <= "111111100111";
      when "001100010011000" => color_data <= "111111111011";
      when "001100010011001" => color_data <= "111111101001";
      when "001100010011010" => color_data <= "111111101010";
      when "001100010011011" => color_data <= "111111101010";
      when "001100010011100" => color_data <= "111111101010";
      when "001100010011101" => color_data <= "111111101010";
      when "001100010011110" => color_data <= "111111101010";
      when "001100010011111" => color_data <= "111111101010";
      when "001100010100000" => color_data <= "111111101010";
      when "001100010100001" => color_data <= "111111101010";
      when "001100010100010" => color_data <= "111111101010";
      when "001100010100011" => color_data <= "111111101010";
      when "001100010100100" => color_data <= "111111101010";
      when "001100010100101" => color_data <= "111111101010";
      when "001100010100110" => color_data <= "111111101010";
      when "001100010100111" => color_data <= "111111101001";
      when "001100010101000" => color_data <= "111111101001";
      when "001100010101001" => color_data <= "111111111011";
      when "001100010101010" => color_data <= "111111010100";
      when "001100010101011" => color_data <= "111111010000";
      when "001100010101100" => color_data <= "111111010000";
      when "001100010101101" => color_data <= "111111010000";
      when "001100010101110" => color_data <= "111111010000";
      when "001100010101111" => color_data <= "111111010000";
      when "001100010110000" => color_data <= "111111010000";
      when "001100010110001" => color_data <= "111111010000";
      when "001100010110010" => color_data <= "111111010000";
      when "001100010110011" => color_data <= "111111010000";
      when "001100010110100" => color_data <= "111111010000";
      when "001100010110101" => color_data <= "111111010000";
      when "001100010110110" => color_data <= "111111010000";
      when "001100010110111" => color_data <= "111111010000";
      when "001100010111000" => color_data <= "111111010000";
      when "001100010111001" => color_data <= "111111010000";
      when "001100010111010" => color_data <= "111111010000";
      when "001100010111011" => color_data <= "111111010001";
      when "001100010111100" => color_data <= "111111101010";
      when "001100010111101" => color_data <= "111111101010";
      when "001100010111110" => color_data <= "111111101001";
      when "001100010111111" => color_data <= "111111101010";
      when "001100011000000" => color_data <= "111111101010";
      when "001100011000001" => color_data <= "111111101010";
      when "001100011000010" => color_data <= "111111101010";
      when "001100011000011" => color_data <= "111111101010";
      when "001100011000100" => color_data <= "111111101010";
      when "001100011000101" => color_data <= "111111101010";
      when "001100011000110" => color_data <= "111111101010";
      when "001100011000111" => color_data <= "111111101010";
      when "001100011001000" => color_data <= "111111101010";
      when "001100011001001" => color_data <= "111111101001";
      when "001100011001010" => color_data <= "111111101010";
      when "001100011001011" => color_data <= "111111111011";
      when "001100011001100" => color_data <= "111111100111";
      when "001100011001101" => color_data <= "111111100101";
      when "001100011001110" => color_data <= "100001110010";
      when "001100011001111" => color_data <= "000000000000";
      when "001100011010000" => color_data <= "000000000000";
      when "001100011010001" => color_data <= "000000000000";
      when "001100011010010" => color_data <= "000000000000";
      when "001100011010011" => color_data <= "000000000000";
      when "001100011010100" => color_data <= "000000000000";
      when "001100011010101" => color_data <= "000000000000";
      when "001100011010110" => color_data <= "000000000000";
      when "001100011010111" => color_data <= "000000000000";
      when "001100011011000" => color_data <= "110110100000";
      when "001100011011001" => color_data <= "111111000000";
      when "001100011011010" => color_data <= "111110110000";
      when "001100011011011" => color_data <= "011001010011";
      when "001100011011100" => color_data <= "000000000000";
      when "001100011011101" => color_data <= "000000000000";
      when "001100011011110" => color_data <= "000000000000";
      when "001100011011111" => color_data <= "000000000000";
      when "001100011100000" => color_data <= "000000000000";
      when "001100011100001" => color_data <= "000000000000";
      when "001100011100010" => color_data <= "000000000000";
      when "001100011100011" => color_data <= "000000000000";
      when "001100100000000" => color_data <= "000000000000";
      when "001100100000001" => color_data <= "000000000000";
      when "001100100000010" => color_data <= "000000000000";
      when "001100100000011" => color_data <= "000000000000";
      when "001100100000100" => color_data <= "000000000000";
      when "001100100000101" => color_data <= "000000000000";
      when "001100100000110" => color_data <= "000000000000";
      when "001100100000111" => color_data <= "000000000000";
      when "001100100001000" => color_data <= "000000000000";
      when "001100100001001" => color_data <= "000000000000";
      when "001100100001010" => color_data <= "000000000000";
      when "001100100001011" => color_data <= "000000000000";
      when "001100100001100" => color_data <= "100001100010";
      when "001100100001101" => color_data <= "111110110000";
      when "001100100001110" => color_data <= "111111000000";
      when "001100100001111" => color_data <= "101110010001";
      when "001100100010000" => color_data <= "000000000000";
      when "001100100010001" => color_data <= "000000000000";
      when "001100100010010" => color_data <= "000000000000";
      when "001100100010011" => color_data <= "000000000000";
      when "001100100010100" => color_data <= "000000000000";
      when "001100100010101" => color_data <= "000000000000";
      when "001100100010110" => color_data <= "100010000010";
      when "001100100010111" => color_data <= "111111100110";
      when "001100100011000" => color_data <= "111111101010";
      when "001100100011001" => color_data <= "111111101010";
      when "001100100011010" => color_data <= "111111101010";
      when "001100100011011" => color_data <= "111111101010";
      when "001100100011100" => color_data <= "111111101010";
      when "001100100011101" => color_data <= "111111101010";
      when "001100100011110" => color_data <= "111111101010";
      when "001100100011111" => color_data <= "111111101010";
      when "001100100100000" => color_data <= "111111101010";
      when "001100100100001" => color_data <= "111111101010";
      when "001100100100010" => color_data <= "111111101010";
      when "001100100100011" => color_data <= "111111101010";
      when "001100100100100" => color_data <= "111111101010";
      when "001100100100101" => color_data <= "111111101010";
      when "001100100100110" => color_data <= "111111101010";
      when "001100100100111" => color_data <= "111111101010";
      when "001100100101000" => color_data <= "111111101001";
      when "001100100101001" => color_data <= "111111111011";
      when "001100100101010" => color_data <= "111111100110";
      when "001100100101011" => color_data <= "111111010000";
      when "001100100101100" => color_data <= "111111010000";
      when "001100100101101" => color_data <= "111111010000";
      when "001100100101110" => color_data <= "111111010000";
      when "001100100101111" => color_data <= "111111010000";
      when "001100100110000" => color_data <= "111111010000";
      when "001100100110001" => color_data <= "111111010000";
      when "001100100110010" => color_data <= "111111010000";
      when "001100100110011" => color_data <= "111111010000";
      when "001100100110100" => color_data <= "111111010000";
      when "001100100110101" => color_data <= "111111010000";
      when "001100100110110" => color_data <= "111111010000";
      when "001100100110111" => color_data <= "111111010000";
      when "001100100111000" => color_data <= "111111010000";
      when "001100100111001" => color_data <= "111111010001";
      when "001100100111010" => color_data <= "111111000000";
      when "001100100111011" => color_data <= "111111010100";
      when "001100100111100" => color_data <= "111111111011";
      when "001100100111101" => color_data <= "111111101001";
      when "001100100111110" => color_data <= "111111101010";
      when "001100100111111" => color_data <= "111111101010";
      when "001100101000000" => color_data <= "111111101010";
      when "001100101000001" => color_data <= "111111101010";
      when "001100101000010" => color_data <= "111111101010";
      when "001100101000011" => color_data <= "111111101010";
      when "001100101000100" => color_data <= "111111101010";
      when "001100101000101" => color_data <= "111111101010";
      when "001100101000110" => color_data <= "111111101010";
      when "001100101000111" => color_data <= "111111101010";
      when "001100101001000" => color_data <= "111111101010";
      when "001100101001001" => color_data <= "111111101010";
      when "001100101001010" => color_data <= "111111101010";
      when "001100101001011" => color_data <= "111111101010";
      when "001100101001100" => color_data <= "111111100110";
      when "001100101001101" => color_data <= "111111010011";
      when "001100101001110" => color_data <= "010101010011";
      when "001100101001111" => color_data <= "000000000000";
      when "001100101010000" => color_data <= "000000000000";
      when "001100101010001" => color_data <= "000000000000";
      when "001100101010010" => color_data <= "000000000000";
      when "001100101010011" => color_data <= "000000000000";
      when "001100101010100" => color_data <= "000000000000";
      when "001100101010101" => color_data <= "000000000000";
      when "001100101010110" => color_data <= "000000000000";
      when "001100101010111" => color_data <= "010101010011";
      when "001100101011000" => color_data <= "110110100000";
      when "001100101011001" => color_data <= "111111000000";
      when "001100101011010" => color_data <= "110110100000";
      when "001100101011011" => color_data <= "000100000000";
      when "001100101011100" => color_data <= "000000000000";
      when "001100101011101" => color_data <= "000000000000";
      when "001100101011110" => color_data <= "000000000000";
      when "001100101011111" => color_data <= "000000000000";
      when "001100101100000" => color_data <= "000000000000";
      when "001100101100001" => color_data <= "000000000000";
      when "001100101100010" => color_data <= "000000000000";
      when "001100101100011" => color_data <= "000000000000";
      when "001100110000000" => color_data <= "000000000000";
      when "001100110000001" => color_data <= "000000000000";
      when "001100110000010" => color_data <= "000000000000";
      when "001100110000011" => color_data <= "000000000000";
      when "001100110000100" => color_data <= "000000000000";
      when "001100110000101" => color_data <= "000000000000";
      when "001100110000110" => color_data <= "000000000000";
      when "001100110000111" => color_data <= "000000000000";
      when "001100110001000" => color_data <= "000000000000";
      when "001100110001001" => color_data <= "000000000000";
      when "001100110001010" => color_data <= "000000000000";
      when "001100110001011" => color_data <= "000000000000";
      when "001100110001100" => color_data <= "000000000000";
      when "001100110001101" => color_data <= "110110100000";
      when "001100110001110" => color_data <= "111111000000";
      when "001100110001111" => color_data <= "110110100000";
      when "001100110010000" => color_data <= "010101010011";
      when "001100110010001" => color_data <= "000000000000";
      when "001100110010010" => color_data <= "000000000000";
      when "001100110010011" => color_data <= "000000000000";
      when "001100110010100" => color_data <= "000000000000";
      when "001100110010101" => color_data <= "000000000000";
      when "001100110010110" => color_data <= "010000110010";
      when "001100110010111" => color_data <= "101010010010";
      when "001100110011000" => color_data <= "111111101001";
      when "001100110011001" => color_data <= "111111111010";
      when "001100110011010" => color_data <= "111111101010";
      when "001100110011011" => color_data <= "111111101010";
      when "001100110011100" => color_data <= "111111101010";
      when "001100110011101" => color_data <= "111111101010";
      when "001100110011110" => color_data <= "111111101010";
      when "001100110011111" => color_data <= "111111101010";
      when "001100110100000" => color_data <= "111111101010";
      when "001100110100001" => color_data <= "111111101010";
      when "001100110100010" => color_data <= "111111101010";
      when "001100110100011" => color_data <= "111111101010";
      when "001100110100100" => color_data <= "111111101010";
      when "001100110100101" => color_data <= "111111101010";
      when "001100110100110" => color_data <= "111111101010";
      when "001100110100111" => color_data <= "111111101010";
      when "001100110101000" => color_data <= "111111101010";
      when "001100110101001" => color_data <= "111111111010";
      when "001100110101010" => color_data <= "111111101001";
      when "001100110101011" => color_data <= "111111010001";
      when "001100110101100" => color_data <= "111111010000";
      when "001100110101101" => color_data <= "111111010000";
      when "001100110101110" => color_data <= "111111010000";
      when "001100110101111" => color_data <= "111111010000";
      when "001100110110000" => color_data <= "111111010000";
      when "001100110110001" => color_data <= "111111010000";
      when "001100110110010" => color_data <= "111111010000";
      when "001100110110011" => color_data <= "111111010000";
      when "001100110110100" => color_data <= "111111010000";
      when "001100110110101" => color_data <= "111111010000";
      when "001100110110110" => color_data <= "111111010000";
      when "001100110110111" => color_data <= "111111010000";
      when "001100110111000" => color_data <= "111111010000";
      when "001100110111001" => color_data <= "111111010000";
      when "001100110111010" => color_data <= "111111010000";
      when "001100110111011" => color_data <= "111111101000";
      when "001100110111100" => color_data <= "111111111011";
      when "001100110111101" => color_data <= "111111101010";
      when "001100110111110" => color_data <= "111111101010";
      when "001100110111111" => color_data <= "111111101010";
      when "001100111000000" => color_data <= "111111101010";
      when "001100111000001" => color_data <= "111111101010";
      when "001100111000010" => color_data <= "111111101010";
      when "001100111000011" => color_data <= "111111101010";
      when "001100111000100" => color_data <= "111111101010";
      when "001100111000101" => color_data <= "111111101010";
      when "001100111000110" => color_data <= "111111101010";
      when "001100111000111" => color_data <= "111111101010";
      when "001100111001000" => color_data <= "111111101010";
      when "001100111001001" => color_data <= "111111101010";
      when "001100111001010" => color_data <= "111111111010";
      when "001100111001011" => color_data <= "111111100111";
      when "001100111001100" => color_data <= "111111100101";
      when "001100111001101" => color_data <= "100001110010";
      when "001100111001110" => color_data <= "000100010001";
      when "001100111001111" => color_data <= "000000000000";
      when "001100111010000" => color_data <= "000000000000";
      when "001100111010001" => color_data <= "000000000000";
      when "001100111010010" => color_data <= "000000000000";
      when "001100111010011" => color_data <= "000000000000";
      when "001100111010100" => color_data <= "000000000000";
      when "001100111010101" => color_data <= "000000000000";
      when "001100111010110" => color_data <= "000000000000";
      when "001100111010111" => color_data <= "110010010001";
      when "001100111011000" => color_data <= "111111000000";
      when "001100111011001" => color_data <= "111110110000";
      when "001100111011010" => color_data <= "100001110010";
      when "001100111011011" => color_data <= "000000000000";
      when "001100111011100" => color_data <= "000000000000";
      when "001100111011101" => color_data <= "000000000000";
      when "001100111011110" => color_data <= "000000000000";
      when "001100111011111" => color_data <= "000000000000";
      when "001100111100000" => color_data <= "000000000000";
      when "001100111100001" => color_data <= "000000000000";
      when "001100111100010" => color_data <= "000000000000";
      when "001100111100011" => color_data <= "000000000000";
      when "001101000000000" => color_data <= "000000000000";
      when "001101000000001" => color_data <= "000000000000";
      when "001101000000010" => color_data <= "000000000000";
      when "001101000000011" => color_data <= "000000000000";
      when "001101000000100" => color_data <= "000000000000";
      when "001101000000101" => color_data <= "000000000000";
      when "001101000000110" => color_data <= "000000000000";
      when "001101000000111" => color_data <= "000000000000";
      when "001101000001000" => color_data <= "000000000000";
      when "001101000001001" => color_data <= "000000000000";
      when "001101000001010" => color_data <= "000000000000";
      when "001101000001011" => color_data <= "000000000000";
      when "001101000001100" => color_data <= "000000000000";
      when "001101000001101" => color_data <= "100001110010";
      when "001101000001110" => color_data <= "111110110000";
      when "001101000001111" => color_data <= "111111000000";
      when "001101000010000" => color_data <= "110010010000";
      when "001101000010001" => color_data <= "000000000000";
      when "001101000010010" => color_data <= "000000000000";
      when "001101000010011" => color_data <= "000000000000";
      when "001101000010100" => color_data <= "000000000000";
      when "001101000010101" => color_data <= "000000000000";
      when "001101000010110" => color_data <= "000000000000";
      when "001101000010111" => color_data <= "101010010010";
      when "001101000011000" => color_data <= "111111100110";
      when "001101000011001" => color_data <= "111111111011";
      when "001101000011010" => color_data <= "111111101001";
      when "001101000011011" => color_data <= "111111101010";
      when "001101000011100" => color_data <= "111111101010";
      when "001101000011101" => color_data <= "111111101010";
      when "001101000011110" => color_data <= "111111101010";
      when "001101000011111" => color_data <= "111111101010";
      when "001101000100000" => color_data <= "111111101010";
      when "001101000100001" => color_data <= "111111101010";
      when "001101000100010" => color_data <= "111111101010";
      when "001101000100011" => color_data <= "111111101010";
      when "001101000100100" => color_data <= "111111101010";
      when "001101000100101" => color_data <= "111111101010";
      when "001101000100110" => color_data <= "111111101010";
      when "001101000100111" => color_data <= "111111101010";
      when "001101000101000" => color_data <= "111111101010";
      when "001101000101001" => color_data <= "111111101010";
      when "001101000101010" => color_data <= "111111111011";
      when "001101000101011" => color_data <= "111111100101";
      when "001101000101100" => color_data <= "111111000000";
      when "001101000101101" => color_data <= "111111010000";
      when "001101000101110" => color_data <= "111111010000";
      when "001101000101111" => color_data <= "111111010000";
      when "001101000110000" => color_data <= "111111010000";
      when "001101000110001" => color_data <= "111111010000";
      when "001101000110010" => color_data <= "111111010000";
      when "001101000110011" => color_data <= "111111010000";
      when "001101000110100" => color_data <= "111111010000";
      when "001101000110101" => color_data <= "111111010000";
      when "001101000110110" => color_data <= "111111010000";
      when "001101000110111" => color_data <= "111111010000";
      when "001101000111000" => color_data <= "111111010000";
      when "001101000111001" => color_data <= "111111000000";
      when "001101000111010" => color_data <= "111111010011";
      when "001101000111011" => color_data <= "111111111011";
      when "001101000111100" => color_data <= "111111101001";
      when "001101000111101" => color_data <= "111111101010";
      when "001101000111110" => color_data <= "111111101010";
      when "001101000111111" => color_data <= "111111101010";
      when "001101001000000" => color_data <= "111111101010";
      when "001101001000001" => color_data <= "111111101010";
      when "001101001000010" => color_data <= "111111101010";
      when "001101001000011" => color_data <= "111111101010";
      when "001101001000100" => color_data <= "111111101010";
      when "001101001000101" => color_data <= "111111101010";
      when "001101001000110" => color_data <= "111111101010";
      when "001101001000111" => color_data <= "111111101010";
      when "001101001001000" => color_data <= "111111101010";
      when "001101001001001" => color_data <= "111111101001";
      when "001101001001010" => color_data <= "111111111011";
      when "001101001001011" => color_data <= "111111100110";
      when "001101001001100" => color_data <= "111111010100";
      when "001101001001101" => color_data <= "011001010011";
      when "001101001001110" => color_data <= "000000000000";
      when "001101001001111" => color_data <= "000000000000";
      when "001101001010000" => color_data <= "000000000000";
      when "001101001010001" => color_data <= "000000000000";
      when "001101001010010" => color_data <= "000000000000";
      when "001101001010011" => color_data <= "000000000000";
      when "001101001010100" => color_data <= "000000000000";
      when "001101001010101" => color_data <= "000000000000";
      when "001101001010110" => color_data <= "010101000010";
      when "001101001010111" => color_data <= "110110100000";
      when "001101001011000" => color_data <= "111111000000";
      when "001101001011001" => color_data <= "110110100000";
      when "001101001011010" => color_data <= "000100000000";
      when "001101001011011" => color_data <= "000000000000";
      when "001101001011100" => color_data <= "000000000000";
      when "001101001011101" => color_data <= "000000000000";
      when "001101001011110" => color_data <= "000000000000";
      when "001101001011111" => color_data <= "000000000000";
      when "001101001100000" => color_data <= "000000000000";
      when "001101001100001" => color_data <= "000000000000";
      when "001101001100010" => color_data <= "000000000000";
      when "001101001100011" => color_data <= "000000000000";
      when "001101010000000" => color_data <= "000000000000";
      when "001101010000001" => color_data <= "000000000000";
      when "001101010000010" => color_data <= "000000000000";
      when "001101010000011" => color_data <= "000000000000";
      when "001101010000100" => color_data <= "000000000000";
      when "001101010000101" => color_data <= "000000000000";
      when "001101010000110" => color_data <= "000000000000";
      when "001101010000111" => color_data <= "000000000000";
      when "001101010001000" => color_data <= "000000000000";
      when "001101010001001" => color_data <= "000000000000";
      when "001101010001010" => color_data <= "000000000000";
      when "001101010001011" => color_data <= "000000000000";
      when "001101010001100" => color_data <= "000000000000";
      when "001101010001101" => color_data <= "000100010001";
      when "001101010001110" => color_data <= "110110100000";
      when "001101010001111" => color_data <= "111111000001";
      when "001101010010000" => color_data <= "110110100000";
      when "001101010010001" => color_data <= "011001010011";
      when "001101010010010" => color_data <= "000000000000";
      when "001101010010011" => color_data <= "000000000000";
      when "001101010010100" => color_data <= "000000000000";
      when "001101010010101" => color_data <= "000000000000";
      when "001101010010110" => color_data <= "000000000000";
      when "001101010010111" => color_data <= "010101000010";
      when "001101010011000" => color_data <= "101010010010";
      when "001101010011001" => color_data <= "111111111010";
      when "001101010011010" => color_data <= "111111101010";
      when "001101010011011" => color_data <= "111111101010";
      when "001101010011100" => color_data <= "111111101010";
      when "001101010011101" => color_data <= "111111101010";
      when "001101010011110" => color_data <= "111111101010";
      when "001101010011111" => color_data <= "111111101010";
      when "001101010100000" => color_data <= "111111101010";
      when "001101010100001" => color_data <= "111111101010";
      when "001101010100010" => color_data <= "111111101010";
      when "001101010100011" => color_data <= "111111101010";
      when "001101010100100" => color_data <= "111111101010";
      when "001101010100101" => color_data <= "111111101010";
      when "001101010100110" => color_data <= "111111101010";
      when "001101010100111" => color_data <= "111111101010";
      when "001101010101000" => color_data <= "111111101001";
      when "001101010101001" => color_data <= "111111101001";
      when "001101010101010" => color_data <= "111111111011";
      when "001101010101011" => color_data <= "111111101000";
      when "001101010101100" => color_data <= "111111010010";
      when "001101010101101" => color_data <= "111111010010";
      when "001101010101110" => color_data <= "111111010001";
      when "001101010101111" => color_data <= "111111010001";
      when "001101010110000" => color_data <= "111111010001";
      when "001101010110001" => color_data <= "111111010001";
      when "001101010110010" => color_data <= "111111010001";
      when "001101010110011" => color_data <= "111111010001";
      when "001101010110100" => color_data <= "111111010001";
      when "001101010110101" => color_data <= "111111010001";
      when "001101010110110" => color_data <= "111111010001";
      when "001101010110111" => color_data <= "111111010001";
      when "001101010111000" => color_data <= "111111010010";
      when "001101010111001" => color_data <= "111111010010";
      when "001101010111010" => color_data <= "111111100110";
      when "001101010111011" => color_data <= "111111111011";
      when "001101010111100" => color_data <= "111111101001";
      when "001101010111101" => color_data <= "111111101010";
      when "001101010111110" => color_data <= "111111101010";
      when "001101010111111" => color_data <= "111111101010";
      when "001101011000000" => color_data <= "111111101010";
      when "001101011000001" => color_data <= "111111101010";
      when "001101011000010" => color_data <= "111111101010";
      when "001101011000011" => color_data <= "111111101010";
      when "001101011000100" => color_data <= "111111101010";
      when "001101011000101" => color_data <= "111111101010";
      when "001101011000110" => color_data <= "111111101010";
      when "001101011000111" => color_data <= "111111101010";
      when "001101011001000" => color_data <= "111111101010";
      when "001101011001001" => color_data <= "111111111011";
      when "001101011001010" => color_data <= "111111101000";
      when "001101011001011" => color_data <= "111111100101";
      when "001101011001100" => color_data <= "100110000010";
      when "001101011001101" => color_data <= "001000100001";
      when "001101011001110" => color_data <= "000000000000";
      when "001101011001111" => color_data <= "000000000000";
      when "001101011010000" => color_data <= "000000000000";
      when "001101011010001" => color_data <= "000000000000";
      when "001101011010010" => color_data <= "000000000000";
      when "001101011010011" => color_data <= "000000000000";
      when "001101011010100" => color_data <= "000000000000";
      when "001101011010101" => color_data <= "000000000000";
      when "001101011010110" => color_data <= "110010010001";
      when "001101011010111" => color_data <= "111111000000";
      when "001101011011000" => color_data <= "111110110000";
      when "001101011011001" => color_data <= "100101110010";
      when "001101011011010" => color_data <= "000000000000";
      when "001101011011011" => color_data <= "000000000000";
      when "001101011011100" => color_data <= "000000000000";
      when "001101011011101" => color_data <= "000000000000";
      when "001101011011110" => color_data <= "000000000000";
      when "001101011011111" => color_data <= "000000000000";
      when "001101011100000" => color_data <= "000000000000";
      when "001101011100001" => color_data <= "000000000000";
      when "001101011100010" => color_data <= "000000000000";
      when "001101011100011" => color_data <= "000000000000";
      when "001101100000000" => color_data <= "000000000000";
      when "001101100000001" => color_data <= "000000000000";
      when "001101100000010" => color_data <= "000000000000";
      when "001101100000011" => color_data <= "000000000000";
      when "001101100000100" => color_data <= "000000000000";
      when "001101100000101" => color_data <= "000000000000";
      when "001101100000110" => color_data <= "000000000000";
      when "001101100000111" => color_data <= "000000000000";
      when "001101100001000" => color_data <= "000000000000";
      when "001101100001001" => color_data <= "000000000000";
      when "001101100001010" => color_data <= "000000000000";
      when "001101100001011" => color_data <= "000000000000";
      when "001101100001100" => color_data <= "000000000000";
      when "001101100001101" => color_data <= "000000000000";
      when "001101100001110" => color_data <= "100110000010";
      when "001101100001111" => color_data <= "111110110000";
      when "001101100010000" => color_data <= "111111000000";
      when "001101100010001" => color_data <= "110010010001";
      when "001101100010010" => color_data <= "000000000000";
      when "001101100010011" => color_data <= "000000000000";
      when "001101100010100" => color_data <= "000000000000";
      when "001101100010101" => color_data <= "000000000000";
      when "001101100010110" => color_data <= "000000000000";
      when "001101100010111" => color_data <= "000000000000";
      when "001101100011000" => color_data <= "101010010010";
      when "001101100011001" => color_data <= "111111100111";
      when "001101100011010" => color_data <= "111111111011";
      when "001101100011011" => color_data <= "111111101001";
      when "001101100011100" => color_data <= "111111101010";
      when "001101100011101" => color_data <= "111111101001";
      when "001101100011110" => color_data <= "111111101010";
      when "001101100011111" => color_data <= "111111101010";
      when "001101100100000" => color_data <= "111111101010";
      when "001101100100001" => color_data <= "111111101010";
      when "001101100100010" => color_data <= "111111101010";
      when "001101100100011" => color_data <= "111111101010";
      when "001101100100100" => color_data <= "111111101010";
      when "001101100100101" => color_data <= "111111101010";
      when "001101100100110" => color_data <= "111111101010";
      when "001101100100111" => color_data <= "111111101001";
      when "001101100101000" => color_data <= "111111101001";
      when "001101100101001" => color_data <= "111111111011";
      when "001101100101010" => color_data <= "111111101001";
      when "001101100101011" => color_data <= "111111100101";
      when "001101100101100" => color_data <= "111111100111";
      when "001101100101101" => color_data <= "111111100111";
      when "001101100101110" => color_data <= "111111100111";
      when "001101100101111" => color_data <= "111111100110";
      when "001101100110000" => color_data <= "111111100110";
      when "001101100110001" => color_data <= "111111100110";
      when "001101100110010" => color_data <= "111111100110";
      when "001101100110011" => color_data <= "111111100110";
      when "001101100110100" => color_data <= "111111100110";
      when "001101100110101" => color_data <= "111111100110";
      when "001101100110110" => color_data <= "111111100110";
      when "001101100110111" => color_data <= "111111100110";
      when "001101100111000" => color_data <= "111111100111";
      when "001101100111001" => color_data <= "111111101000";
      when "001101100111010" => color_data <= "111111100101";
      when "001101100111011" => color_data <= "111111101000";
      when "001101100111100" => color_data <= "111111101011";
      when "001101100111101" => color_data <= "111111101010";
      when "001101100111110" => color_data <= "111111101010";
      when "001101100111111" => color_data <= "111111101010";
      when "001101101000000" => color_data <= "111111101010";
      when "001101101000001" => color_data <= "111111101010";
      when "001101101000010" => color_data <= "111111101010";
      when "001101101000011" => color_data <= "111111101010";
      when "001101101000100" => color_data <= "111111101010";
      when "001101101000101" => color_data <= "111111101010";
      when "001101101000110" => color_data <= "111111101010";
      when "001101101000111" => color_data <= "111111101001";
      when "001101101001000" => color_data <= "111111101010";
      when "001101101001001" => color_data <= "111111111010";
      when "001101101001010" => color_data <= "111111100110";
      when "001101101001011" => color_data <= "111111010100";
      when "001101101001100" => color_data <= "011001100011";
      when "001101101001101" => color_data <= "000000000000";
      when "001101101001110" => color_data <= "000000000000";
      when "001101101001111" => color_data <= "000000000000";
      when "001101101010000" => color_data <= "000000000000";
      when "001101101010001" => color_data <= "000000000000";
      when "001101101010010" => color_data <= "000000000000";
      when "001101101010011" => color_data <= "000000000000";
      when "001101101010100" => color_data <= "000000000000";
      when "001101101010101" => color_data <= "010101000010";
      when "001101101010110" => color_data <= "110110100000";
      when "001101101010111" => color_data <= "111111000001";
      when "001101101011000" => color_data <= "110110100000";
      when "001101101011001" => color_data <= "001000100001";
      when "001101101011010" => color_data <= "000000000000";
      when "001101101011011" => color_data <= "000000000000";
      when "001101101011100" => color_data <= "000000000000";
      when "001101101011101" => color_data <= "000000000000";
      when "001101101011110" => color_data <= "000000000000";
      when "001101101011111" => color_data <= "000000000000";
      when "001101101100000" => color_data <= "000000000000";
      when "001101101100001" => color_data <= "000000000000";
      when "001101101100010" => color_data <= "000000000000";
      when "001101101100011" => color_data <= "000000000000";
      when "001101110000000" => color_data <= "000000000000";
      when "001101110000001" => color_data <= "000000000000";
      when "001101110000010" => color_data <= "000000000000";
      when "001101110000011" => color_data <= "000000000000";
      when "001101110000100" => color_data <= "000000000000";
      when "001101110000101" => color_data <= "000000000000";
      when "001101110000110" => color_data <= "000000000000";
      when "001101110000111" => color_data <= "000000000000";
      when "001101110001000" => color_data <= "000000000000";
      when "001101110001001" => color_data <= "000000000000";
      when "001101110001010" => color_data <= "000000000000";
      when "001101110001011" => color_data <= "000000000000";
      when "001101110001100" => color_data <= "000000000000";
      when "001101110001101" => color_data <= "000000000000";
      when "001101110001110" => color_data <= "000100010001";
      when "001101110001111" => color_data <= "110110100000";
      when "001101110010000" => color_data <= "111111000000";
      when "001101110010001" => color_data <= "110110100000";
      when "001101110010010" => color_data <= "011001100011";
      when "001101110010011" => color_data <= "000000000000";
      when "001101110010100" => color_data <= "000000000000";
      when "001101110010101" => color_data <= "000000000000";
      when "001101110010110" => color_data <= "000000000000";
      when "001101110010111" => color_data <= "000000000000";
      when "001101110011000" => color_data <= "001100110010";
      when "001101110011001" => color_data <= "101110100001";
      when "001101110011010" => color_data <= "111111111010";
      when "001101110011011" => color_data <= "111111111011";
      when "001101110011100" => color_data <= "111111101010";
      when "001101110011101" => color_data <= "111111101010";
      when "001101110011110" => color_data <= "111111101010";
      when "001101110011111" => color_data <= "111111101010";
      when "001101110100000" => color_data <= "111111101010";
      when "001101110100001" => color_data <= "111111101010";
      when "001101110100010" => color_data <= "111111101010";
      when "001101110100011" => color_data <= "111111101010";
      when "001101110100100" => color_data <= "111111101010";
      when "001101110100101" => color_data <= "111111101010";
      when "001101110100110" => color_data <= "111111101010";
      when "001101110100111" => color_data <= "111111101001";
      when "001101110101000" => color_data <= "111111111011";
      when "001101110101001" => color_data <= "111111101001";
      when "001101110101010" => color_data <= "111111010100";
      when "001101110101011" => color_data <= "111111100110";
      when "001101110101100" => color_data <= "111111100111";
      when "001101110101101" => color_data <= "111111100111";
      when "001101110101110" => color_data <= "111111100111";
      when "001101110101111" => color_data <= "111111100111";
      when "001101110110000" => color_data <= "111111100111";
      when "001101110110001" => color_data <= "111111100111";
      when "001101110110010" => color_data <= "111111100111";
      when "001101110110011" => color_data <= "111111100111";
      when "001101110110100" => color_data <= "111111100111";
      when "001101110110101" => color_data <= "111111100111";
      when "001101110110110" => color_data <= "111111100111";
      when "001101110110111" => color_data <= "111111100111";
      when "001101110111000" => color_data <= "111111100111";
      when "001101110111001" => color_data <= "111111100111";
      when "001101110111010" => color_data <= "111111100101";
      when "001101110111011" => color_data <= "111111100110";
      when "001101110111100" => color_data <= "111111111010";
      when "001101110111101" => color_data <= "111111101001";
      when "001101110111110" => color_data <= "111111101010";
      when "001101110111111" => color_data <= "111111101010";
      when "001101111000000" => color_data <= "111111101010";
      when "001101111000001" => color_data <= "111111101010";
      when "001101111000010" => color_data <= "111111101010";
      when "001101111000011" => color_data <= "111111101010";
      when "001101111000100" => color_data <= "111111101010";
      when "001101111000101" => color_data <= "111111101010";
      when "001101111000110" => color_data <= "111111101001";
      when "001101111000111" => color_data <= "111111101010";
      when "001101111001000" => color_data <= "111111111100";
      when "001101111001001" => color_data <= "111111100111";
      when "001101111001010" => color_data <= "111111100101";
      when "001101111001011" => color_data <= "100001110010";
      when "001101111001100" => color_data <= "000000000000";
      when "001101111001101" => color_data <= "000000000000";
      when "001101111001110" => color_data <= "000000000000";
      when "001101111001111" => color_data <= "000000000000";
      when "001101111010000" => color_data <= "000000000000";
      when "001101111010001" => color_data <= "000000000000";
      when "001101111010010" => color_data <= "000000000000";
      when "001101111010011" => color_data <= "000000000000";
      when "001101111010100" => color_data <= "000000000000";
      when "001101111010101" => color_data <= "110010100000";
      when "001101111010110" => color_data <= "111111000000";
      when "001101111010111" => color_data <= "111110110000";
      when "001101111011000" => color_data <= "100110000010";
      when "001101111011001" => color_data <= "000000000000";
      when "001101111011010" => color_data <= "000000000000";
      when "001101111011011" => color_data <= "000000000000";
      when "001101111011100" => color_data <= "000000000000";
      when "001101111011101" => color_data <= "000000000000";
      when "001101111011110" => color_data <= "000000000000";
      when "001101111011111" => color_data <= "000000000000";
      when "001101111100000" => color_data <= "000000000000";
      when "001101111100001" => color_data <= "000000000000";
      when "001101111100010" => color_data <= "000000000000";
      when "001101111100011" => color_data <= "000000000000";
      when "001110000000000" => color_data <= "000000000000";
      when "001110000000001" => color_data <= "000000000000";
      when "001110000000010" => color_data <= "000000000000";
      when "001110000000011" => color_data <= "000000000000";
      when "001110000000100" => color_data <= "000000000000";
      when "001110000000101" => color_data <= "000000000000";
      when "001110000000110" => color_data <= "000000000000";
      when "001110000000111" => color_data <= "000000000000";
      when "001110000001000" => color_data <= "000000000000";
      when "001110000001001" => color_data <= "000000000000";
      when "001110000001010" => color_data <= "000000000000";
      when "001110000001011" => color_data <= "000000000000";
      when "001110000001100" => color_data <= "000000000000";
      when "001110000001101" => color_data <= "000000000000";
      when "001110000001110" => color_data <= "000000000000";
      when "001110000001111" => color_data <= "100001110010";
      when "001110000010000" => color_data <= "111110110000";
      when "001110000010001" => color_data <= "111111000000";
      when "001110000010010" => color_data <= "110110100000";
      when "001110000010011" => color_data <= "000000000000";
      when "001110000010100" => color_data <= "000000000000";
      when "001110000010101" => color_data <= "000000000000";
      when "001110000010110" => color_data <= "000000000000";
      when "001110000010111" => color_data <= "000000000000";
      when "001110000011000" => color_data <= "000000000000";
      when "001110000011001" => color_data <= "100110000010";
      when "001110000011010" => color_data <= "110110110000";
      when "001110000011011" => color_data <= "111111101000";
      when "001110000011100" => color_data <= "111111111011";
      when "001110000011101" => color_data <= "111111111011";
      when "001110000011110" => color_data <= "111111111010";
      when "001110000011111" => color_data <= "111111101001";
      when "001110000100000" => color_data <= "111111101010";
      when "001110000100001" => color_data <= "111111101010";
      when "001110000100010" => color_data <= "111111101010";
      when "001110000100011" => color_data <= "111111101010";
      when "001110000100100" => color_data <= "111111101010";
      when "001110000100101" => color_data <= "111111101010";
      when "001110000100110" => color_data <= "111111101010";
      when "001110000100111" => color_data <= "111111111011";
      when "001110000101000" => color_data <= "111111101000";
      when "001110000101001" => color_data <= "111111010100";
      when "001110000101010" => color_data <= "111111100110";
      when "001110000101011" => color_data <= "111111100111";
      when "001110000101100" => color_data <= "111111100111";
      when "001110000101101" => color_data <= "111111100111";
      when "001110000101110" => color_data <= "111111100111";
      when "001110000101111" => color_data <= "111111100111";
      when "001110000110000" => color_data <= "111111100111";
      when "001110000110001" => color_data <= "111111100111";
      when "001110000110010" => color_data <= "111111100111";
      when "001110000110011" => color_data <= "111111100111";
      when "001110000110100" => color_data <= "111111100111";
      when "001110000110101" => color_data <= "111111100111";
      when "001110000110110" => color_data <= "111111100111";
      when "001110000110111" => color_data <= "111111100111";
      when "001110000111000" => color_data <= "111111100111";
      when "001110000111001" => color_data <= "111111100110";
      when "001110000111010" => color_data <= "111111100111";
      when "001110000111011" => color_data <= "111111100101";
      when "001110000111100" => color_data <= "111111101000";
      when "001110000111101" => color_data <= "111111111010";
      when "001110000111110" => color_data <= "111111101001";
      when "001110000111111" => color_data <= "111111101010";
      when "001110001000000" => color_data <= "111111101010";
      when "001110001000001" => color_data <= "111111101010";
      when "001110001000010" => color_data <= "111111101010";
      when "001110001000011" => color_data <= "111111101010";
      when "001110001000100" => color_data <= "111111101001";
      when "001110001000101" => color_data <= "111111101010";
      when "001110001000110" => color_data <= "111111111011";
      when "001110001000111" => color_data <= "111111111010";
      when "001110001001000" => color_data <= "111111010101";
      when "001110001001001" => color_data <= "111111010000";
      when "001110001001010" => color_data <= "101110100001";
      when "001110001001011" => color_data <= "001100110010";
      when "001110001001100" => color_data <= "000000000000";
      when "001110001001101" => color_data <= "000000000000";
      when "001110001001110" => color_data <= "000000000000";
      when "001110001001111" => color_data <= "000000000000";
      when "001110001010000" => color_data <= "000000000000";
      when "001110001010001" => color_data <= "000000000000";
      when "001110001010010" => color_data <= "000000000000";
      when "001110001010011" => color_data <= "000000000000";
      when "001110001010100" => color_data <= "011001100011";
      when "001110001010101" => color_data <= "110110100000";
      when "001110001010110" => color_data <= "111111000000";
      when "001110001010111" => color_data <= "110110100000";
      when "001110001011000" => color_data <= "000100010001";
      when "001110001011001" => color_data <= "000000000000";
      when "001110001011010" => color_data <= "000000000000";
      when "001110001011011" => color_data <= "000000000000";
      when "001110001011100" => color_data <= "000000000000";
      when "001110001011101" => color_data <= "000000000000";
      when "001110001011110" => color_data <= "000000000000";
      when "001110001011111" => color_data <= "000000000000";
      when "001110001100000" => color_data <= "000000000000";
      when "001110001100001" => color_data <= "000000000000";
      when "001110001100010" => color_data <= "000000000000";
      when "001110001100011" => color_data <= "000000000000";
      when "001110010000000" => color_data <= "000000000000";
      when "001110010000001" => color_data <= "000000000000";
      when "001110010000010" => color_data <= "000000000000";
      when "001110010000011" => color_data <= "000000000000";
      when "001110010000100" => color_data <= "000000000000";
      when "001110010000101" => color_data <= "000000000000";
      when "001110010000110" => color_data <= "000000000000";
      when "001110010000111" => color_data <= "000000000000";
      when "001110010001000" => color_data <= "000000000000";
      when "001110010001001" => color_data <= "000000000000";
      when "001110010001010" => color_data <= "000000000000";
      when "001110010001011" => color_data <= "000000000000";
      when "001110010001100" => color_data <= "000000000000";
      when "001110010001101" => color_data <= "000000000000";
      when "001110010001110" => color_data <= "000000000000";
      when "001110010001111" => color_data <= "000100010001";
      when "001110010010000" => color_data <= "110110100000";
      when "001110010010001" => color_data <= "111111000001";
      when "001110010010010" => color_data <= "111110110000";
      when "001110010010011" => color_data <= "100001110010";
      when "001110010010100" => color_data <= "000000000000";
      when "001110010010101" => color_data <= "000000000000";
      when "001110010010110" => color_data <= "000000000000";
      when "001110010010111" => color_data <= "000000000000";
      when "001110010011000" => color_data <= "000000000000";
      when "001110010011001" => color_data <= "000000000000";
      when "001110010011010" => color_data <= "110110110000";
      when "001110010011011" => color_data <= "111111000000";
      when "001110010011100" => color_data <= "111111010011";
      when "001110010011101" => color_data <= "111111100110";
      when "001110010011110" => color_data <= "111111101010";
      when "001110010011111" => color_data <= "111111111011";
      when "001110010100000" => color_data <= "111111111010";
      when "001110010100001" => color_data <= "111111101010";
      when "001110010100010" => color_data <= "111111101010";
      when "001110010100011" => color_data <= "111111101010";
      when "001110010100100" => color_data <= "111111101001";
      when "001110010100101" => color_data <= "111111101001";
      when "001110010100110" => color_data <= "111111111011";
      when "001110010100111" => color_data <= "111111100111";
      when "001110010101000" => color_data <= "111111010100";
      when "001110010101001" => color_data <= "111111100110";
      when "001110010101010" => color_data <= "111111100111";
      when "001110010101011" => color_data <= "111111100111";
      when "001110010101100" => color_data <= "111111100111";
      when "001110010101101" => color_data <= "111111100111";
      when "001110010101110" => color_data <= "111111100111";
      when "001110010101111" => color_data <= "111111100111";
      when "001110010110000" => color_data <= "111111100111";
      when "001110010110001" => color_data <= "111111100111";
      when "001110010110010" => color_data <= "111111100111";
      when "001110010110011" => color_data <= "111111100111";
      when "001110010110100" => color_data <= "111111100111";
      when "001110010110101" => color_data <= "111111100111";
      when "001110010110110" => color_data <= "111111100111";
      when "001110010110111" => color_data <= "111111100111";
      when "001110010111000" => color_data <= "111111100111";
      when "001110010111001" => color_data <= "111111100111";
      when "001110010111010" => color_data <= "111111100111";
      when "001110010111011" => color_data <= "111111100110";
      when "001110010111100" => color_data <= "111111100101";
      when "001110010111101" => color_data <= "111111111010";
      when "001110010111110" => color_data <= "111111101010";
      when "001110010111111" => color_data <= "111111101010";
      when "001110011000000" => color_data <= "111111101010";
      when "001110011000001" => color_data <= "111111101010";
      when "001110011000010" => color_data <= "111111101001";
      when "001110011000011" => color_data <= "111111101010";
      when "001110011000100" => color_data <= "111111111011";
      when "001110011000101" => color_data <= "111111111011";
      when "001110011000110" => color_data <= "111111100110";
      when "001110011000111" => color_data <= "111111010010";
      when "001110011001000" => color_data <= "111111010000";
      when "001110011001001" => color_data <= "110110110000";
      when "001110011001010" => color_data <= "100001110010";
      when "001110011001011" => color_data <= "000000000000";
      when "001110011001100" => color_data <= "000000000000";
      when "001110011001101" => color_data <= "000000000000";
      when "001110011001110" => color_data <= "000000000000";
      when "001110011001111" => color_data <= "000000000000";
      when "001110011010000" => color_data <= "000000000000";
      when "001110011010001" => color_data <= "000000000000";
      when "001110011010010" => color_data <= "000000000000";
      when "001110011010011" => color_data <= "000000000000";
      when "001110011010100" => color_data <= "110110100000";
      when "001110011010101" => color_data <= "111111000000";
      when "001110011010110" => color_data <= "111110110000";
      when "001110011010111" => color_data <= "100110000010";
      when "001110011011000" => color_data <= "000000000000";
      when "001110011011001" => color_data <= "000000000000";
      when "001110011011010" => color_data <= "000000000000";
      when "001110011011011" => color_data <= "000000000000";
      when "001110011011100" => color_data <= "000000000000";
      when "001110011011101" => color_data <= "000000000000";
      when "001110011011110" => color_data <= "000000000000";
      when "001110011011111" => color_data <= "000000000000";
      when "001110011100000" => color_data <= "000000000000";
      when "001110011100001" => color_data <= "000000000000";
      when "001110011100010" => color_data <= "000000000000";
      when "001110011100011" => color_data <= "000000000000";
      when "001110100000000" => color_data <= "000000000000";
      when "001110100000001" => color_data <= "000000000000";
      when "001110100000010" => color_data <= "000000000000";
      when "001110100000011" => color_data <= "000000000000";
      when "001110100000100" => color_data <= "000000000000";
      when "001110100000101" => color_data <= "000000000000";
      when "001110100000110" => color_data <= "000000000000";
      when "001110100000111" => color_data <= "000000000000";
      when "001110100001000" => color_data <= "000000000000";
      when "001110100001001" => color_data <= "000000000000";
      when "001110100001010" => color_data <= "000000000000";
      when "001110100001011" => color_data <= "000000000000";
      when "001110100001100" => color_data <= "000000000000";
      when "001110100001101" => color_data <= "000000000000";
      when "001110100001110" => color_data <= "000000000000";
      when "001110100001111" => color_data <= "000000000000";
      when "001110100010000" => color_data <= "100001110010";
      when "001110100010001" => color_data <= "111110110000";
      when "001110100010010" => color_data <= "111111000000";
      when "001110100010011" => color_data <= "110110100000";
      when "001110100010100" => color_data <= "000100010001";
      when "001110100010101" => color_data <= "000000000000";
      when "001110100010110" => color_data <= "000000000000";
      when "001110100010111" => color_data <= "000000000000";
      when "001110100011000" => color_data <= "000000000000";
      when "001110100011001" => color_data <= "000000000000";
      when "001110100011010" => color_data <= "000000000000";
      when "001110100011011" => color_data <= "110110110000";
      when "001110100011100" => color_data <= "111111000000";
      when "001110100011101" => color_data <= "111111000000";
      when "001110100011110" => color_data <= "111111010001";
      when "001110100011111" => color_data <= "111111100101";
      when "001110100100000" => color_data <= "111111101001";
      when "001110100100001" => color_data <= "111111101010";
      when "001110100100010" => color_data <= "111111111011";
      when "001110100100011" => color_data <= "111111111011";
      when "001110100100100" => color_data <= "111111111010";
      when "001110100100101" => color_data <= "111111111011";
      when "001110100100110" => color_data <= "111111100110";
      when "001110100100111" => color_data <= "111111010100";
      when "001110100101000" => color_data <= "111111100111";
      when "001110100101001" => color_data <= "111111100111";
      when "001110100101010" => color_data <= "111111100111";
      when "001110100101011" => color_data <= "111111100111";
      when "001110100101100" => color_data <= "111111100111";
      when "001110100101101" => color_data <= "111111100111";
      when "001110100101110" => color_data <= "111111100111";
      when "001110100101111" => color_data <= "111111100111";
      when "001110100110000" => color_data <= "111111100111";
      when "001110100110001" => color_data <= "111111100111";
      when "001110100110010" => color_data <= "111111100111";
      when "001110100110011" => color_data <= "111111100111";
      when "001110100110100" => color_data <= "111111100111";
      when "001110100110101" => color_data <= "111111100111";
      when "001110100110110" => color_data <= "111111100111";
      when "001110100110111" => color_data <= "111111100111";
      when "001110100111000" => color_data <= "111111100111";
      when "001110100111001" => color_data <= "111111100111";
      when "001110100111010" => color_data <= "111111100111";
      when "001110100111011" => color_data <= "111111100111";
      when "001110100111100" => color_data <= "111111010100";
      when "001110100111101" => color_data <= "111111100111";
      when "001110100111110" => color_data <= "111111111011";
      when "001110100111111" => color_data <= "111111101001";
      when "001110101000000" => color_data <= "111111101001";
      when "001110101000001" => color_data <= "111111101010";
      when "001110101000010" => color_data <= "111111111011";
      when "001110101000011" => color_data <= "111111111011";
      when "001110101000100" => color_data <= "111111100111";
      when "001110101000101" => color_data <= "111111010011";
      when "001110101000110" => color_data <= "111111010000";
      when "001110101000111" => color_data <= "111111010000";
      when "001110101001000" => color_data <= "111111000000";
      when "001110101001001" => color_data <= "101110010001";
      when "001110101001010" => color_data <= "000000000000";
      when "001110101001011" => color_data <= "000000000000";
      when "001110101001100" => color_data <= "000000000000";
      when "001110101001101" => color_data <= "000000000000";
      when "001110101001110" => color_data <= "000000000000";
      when "001110101001111" => color_data <= "000000000000";
      when "001110101010000" => color_data <= "000000000000";
      when "001110101010001" => color_data <= "000000000000";
      when "001110101010010" => color_data <= "000000000000";
      when "001110101010011" => color_data <= "100001110010";
      when "001110101010100" => color_data <= "111110110000";
      when "001110101010101" => color_data <= "111111000000";
      when "001110101010110" => color_data <= "110110100000";
      when "001110101010111" => color_data <= "000100010001";
      when "001110101011000" => color_data <= "000000000000";
      when "001110101011001" => color_data <= "000000000000";
      when "001110101011010" => color_data <= "000000000000";
      when "001110101011011" => color_data <= "000000000000";
      when "001110101011100" => color_data <= "000000000000";
      when "001110101011101" => color_data <= "000000000000";
      when "001110101011110" => color_data <= "000000000000";
      when "001110101011111" => color_data <= "000000000000";
      when "001110101100000" => color_data <= "000000000000";
      when "001110101100001" => color_data <= "000000000000";
      when "001110101100010" => color_data <= "000000000000";
      when "001110101100011" => color_data <= "000000000000";
      when "001110110000000" => color_data <= "000000000000";
      when "001110110000001" => color_data <= "000000000000";
      when "001110110000010" => color_data <= "000000000000";
      when "001110110000011" => color_data <= "000000000000";
      when "001110110000100" => color_data <= "000000000000";
      when "001110110000101" => color_data <= "000000000000";
      when "001110110000110" => color_data <= "000000000000";
      when "001110110000111" => color_data <= "000000000000";
      when "001110110001000" => color_data <= "000000000000";
      when "001110110001001" => color_data <= "000000000000";
      when "001110110001010" => color_data <= "000000000000";
      when "001110110001011" => color_data <= "000000000000";
      when "001110110001100" => color_data <= "000000000000";
      when "001110110001101" => color_data <= "000000000000";
      when "001110110001110" => color_data <= "000000000000";
      when "001110110001111" => color_data <= "000000000000";
      when "001110110010000" => color_data <= "000000000000";
      when "001110110010001" => color_data <= "110110100000";
      when "001110110010010" => color_data <= "111111000000";
      when "001110110010011" => color_data <= "111110110000";
      when "001110110010100" => color_data <= "101010000010";
      when "001110110010101" => color_data <= "000000000000";
      when "001110110010110" => color_data <= "000000000000";
      when "001110110010111" => color_data <= "000000000000";
      when "001110110011000" => color_data <= "000000000000";
      when "001110110011001" => color_data <= "000000000000";
      when "001110110011010" => color_data <= "000000000000";
      when "001110110011011" => color_data <= "001000100001";
      when "001110110011100" => color_data <= "110110110000";
      when "001110110011101" => color_data <= "111111010000";
      when "001110110011110" => color_data <= "111111010000";
      when "001110110011111" => color_data <= "111111010000";
      when "001110110100000" => color_data <= "111111100111";
      when "001110110100001" => color_data <= "111111010101";
      when "001110110100010" => color_data <= "111111010100";
      when "001110110100011" => color_data <= "111111100111";
      when "001110110100100" => color_data <= "111111101010";
      when "001110110100101" => color_data <= "111111100111";
      when "001110110100110" => color_data <= "111111100100";
      when "001110110100111" => color_data <= "111111100111";
      when "001110110101000" => color_data <= "111111100111";
      when "001110110101001" => color_data <= "111111100111";
      when "001110110101010" => color_data <= "111111100111";
      when "001110110101011" => color_data <= "111111100111";
      when "001110110101100" => color_data <= "111111100111";
      when "001110110101101" => color_data <= "111111100111";
      when "001110110101110" => color_data <= "111111100111";
      when "001110110101111" => color_data <= "111111100111";
      when "001110110110000" => color_data <= "111111100111";
      when "001110110110001" => color_data <= "111111100111";
      when "001110110110010" => color_data <= "111111100111";
      when "001110110110011" => color_data <= "111111100111";
      when "001110110110100" => color_data <= "111111100111";
      when "001110110110101" => color_data <= "111111100111";
      when "001110110110110" => color_data <= "111111100111";
      when "001110110110111" => color_data <= "111111100111";
      when "001110110111000" => color_data <= "111111100111";
      when "001110110111001" => color_data <= "111111100111";
      when "001110110111010" => color_data <= "111111100111";
      when "001110110111011" => color_data <= "111111100111";
      when "001110110111100" => color_data <= "111111100110";
      when "001110110111101" => color_data <= "111111100100";
      when "001110110111110" => color_data <= "111111101001";
      when "001110110111111" => color_data <= "111111111011";
      when "001110111000000" => color_data <= "111111111011";
      when "001110111000001" => color_data <= "111111101010";
      when "001110111000010" => color_data <= "111111100110";
      when "001110111000011" => color_data <= "111111010011";
      when "001110111000100" => color_data <= "111111000000";
      when "001110111000101" => color_data <= "111111010001";
      when "001110111000110" => color_data <= "111111101000";
      when "001110111000111" => color_data <= "111111010000";
      when "001110111001000" => color_data <= "110110110000";
      when "001110111001001" => color_data <= "000000000000";
      when "001110111001010" => color_data <= "000000000000";
      when "001110111001011" => color_data <= "000000000000";
      when "001110111001100" => color_data <= "000000000000";
      when "001110111001101" => color_data <= "000000000000";
      when "001110111001110" => color_data <= "000000000000";
      when "001110111001111" => color_data <= "000000000000";
      when "001110111010000" => color_data <= "000000000000";
      when "001110111010001" => color_data <= "000000000000";
      when "001110111010010" => color_data <= "000100010001";
      when "001110111010011" => color_data <= "110110100000";
      when "001110111010100" => color_data <= "111111000000";
      when "001110111010101" => color_data <= "111110110000";
      when "001110111010110" => color_data <= "100001110010";
      when "001110111010111" => color_data <= "000000000000";
      when "001110111011000" => color_data <= "000000000000";
      when "001110111011001" => color_data <= "000000000000";
      when "001110111011010" => color_data <= "000000000000";
      when "001110111011011" => color_data <= "000000000000";
      when "001110111011100" => color_data <= "000000000000";
      when "001110111011101" => color_data <= "000000000000";
      when "001110111011110" => color_data <= "000000000000";
      when "001110111011111" => color_data <= "000000000000";
      when "001110111100000" => color_data <= "000000000000";
      when "001110111100001" => color_data <= "000000000000";
      when "001110111100010" => color_data <= "000000000000";
      when "001110111100011" => color_data <= "000000000000";
      when "001111000000000" => color_data <= "000000000000";
      when "001111000000001" => color_data <= "000000000000";
      when "001111000000010" => color_data <= "000000000000";
      when "001111000000011" => color_data <= "000000000000";
      when "001111000000100" => color_data <= "000000000000";
      when "001111000000101" => color_data <= "000000000000";
      when "001111000000110" => color_data <= "000000000000";
      when "001111000000111" => color_data <= "000000000000";
      when "001111000001000" => color_data <= "000000000000";
      when "001111000001001" => color_data <= "000000000000";
      when "001111000001010" => color_data <= "000000000000";
      when "001111000001011" => color_data <= "000000000000";
      when "001111000001100" => color_data <= "000000000000";
      when "001111000001101" => color_data <= "000000000000";
      when "001111000001110" => color_data <= "000000000000";
      when "001111000001111" => color_data <= "000000000000";
      when "001111000010000" => color_data <= "000000000000";
      when "001111000010001" => color_data <= "011001100011";
      when "001111000010010" => color_data <= "110110100000";
      when "001111000010011" => color_data <= "111111000001";
      when "001111000010100" => color_data <= "110110100000";
      when "001111000010101" => color_data <= "010000110010";
      when "001111000010110" => color_data <= "000000000000";
      when "001111000010111" => color_data <= "000000000000";
      when "001111000011000" => color_data <= "000000000000";
      when "001111000011001" => color_data <= "000000000000";
      when "001111000011010" => color_data <= "000000000000";
      when "001111000011011" => color_data <= "000000000000";
      when "001111000011100" => color_data <= "010000110010";
      when "001111000011101" => color_data <= "110110110000";
      when "001111000011110" => color_data <= "111111010000";
      when "001111000011111" => color_data <= "111111010010";
      when "001111000100000" => color_data <= "111111101001";
      when "001111000100001" => color_data <= "111111010011";
      when "001111000100010" => color_data <= "111111000000";
      when "001111000100011" => color_data <= "111111010000";
      when "001111000100100" => color_data <= "111111010001";
      when "001111000100101" => color_data <= "111111100101";
      when "001111000100110" => color_data <= "111111101000";
      when "001111000100111" => color_data <= "111111100111";
      when "001111000101000" => color_data <= "111111100111";
      when "001111000101001" => color_data <= "111111100111";
      when "001111000101010" => color_data <= "111111100111";
      when "001111000101011" => color_data <= "111111100111";
      when "001111000101100" => color_data <= "111111100111";
      when "001111000101101" => color_data <= "111111100111";
      when "001111000101110" => color_data <= "111111100111";
      when "001111000101111" => color_data <= "111111100111";
      when "001111000110000" => color_data <= "111111100111";
      when "001111000110001" => color_data <= "111111100111";
      when "001111000110010" => color_data <= "111111100111";
      when "001111000110011" => color_data <= "111111100111";
      when "001111000110100" => color_data <= "111111100111";
      when "001111000110101" => color_data <= "111111100111";
      when "001111000110110" => color_data <= "111111100111";
      when "001111000110111" => color_data <= "111111100111";
      when "001111000111000" => color_data <= "111111100111";
      when "001111000111001" => color_data <= "111111100111";
      when "001111000111010" => color_data <= "111111100111";
      when "001111000111011" => color_data <= "111111100111";
      when "001111000111100" => color_data <= "111111100111";
      when "001111000111101" => color_data <= "111111100101";
      when "001111000111110" => color_data <= "111111100110";
      when "001111000111111" => color_data <= "111111101001";
      when "001111001000000" => color_data <= "111111100101";
      when "001111001000001" => color_data <= "111111010001";
      when "001111001000010" => color_data <= "111111000000";
      when "001111001000011" => color_data <= "111111010000";
      when "001111001000100" => color_data <= "111111010000";
      when "001111001000101" => color_data <= "111111010011";
      when "001111001000110" => color_data <= "011001100011";
      when "001111001000111" => color_data <= "101010000010";
      when "001111001001000" => color_data <= "000100010001";
      when "001111001001001" => color_data <= "000000000000";
      when "001111001001010" => color_data <= "000000000000";
      when "001111001001011" => color_data <= "000000000000";
      when "001111001001100" => color_data <= "000000000000";
      when "001111001001101" => color_data <= "000000000000";
      when "001111001001110" => color_data <= "000000000000";
      when "001111001001111" => color_data <= "000000000000";
      when "001111001010000" => color_data <= "000000000000";
      when "001111001010001" => color_data <= "000000000000";
      when "001111001010010" => color_data <= "101010000010";
      when "001111001010011" => color_data <= "111110110000";
      when "001111001010100" => color_data <= "111111000000";
      when "001111001010101" => color_data <= "110110100000";
      when "001111001010110" => color_data <= "000000000000";
      when "001111001010111" => color_data <= "000000000000";
      when "001111001011000" => color_data <= "000000000000";
      when "001111001011001" => color_data <= "000000000000";
      when "001111001011010" => color_data <= "000000000000";
      when "001111001011011" => color_data <= "000000000000";
      when "001111001011100" => color_data <= "000000000000";
      when "001111001011101" => color_data <= "000000000000";
      when "001111001011110" => color_data <= "000000000000";
      when "001111001011111" => color_data <= "000000000000";
      when "001111001100000" => color_data <= "000000000000";
      when "001111001100001" => color_data <= "000000000000";
      when "001111001100010" => color_data <= "000000000000";
      when "001111001100011" => color_data <= "000000000000";
      when "001111010000000" => color_data <= "000000000000";
      when "001111010000001" => color_data <= "000000000000";
      when "001111010000010" => color_data <= "000000000000";
      when "001111010000011" => color_data <= "000000000000";
      when "001111010000100" => color_data <= "000000000000";
      when "001111010000101" => color_data <= "000000000000";
      when "001111010000110" => color_data <= "000000000000";
      when "001111010000111" => color_data <= "000000000000";
      when "001111010001000" => color_data <= "000000000000";
      when "001111010001001" => color_data <= "000000000000";
      when "001111010001010" => color_data <= "000000000000";
      when "001111010001011" => color_data <= "000000000000";
      when "001111010001100" => color_data <= "000000000000";
      when "001111010001101" => color_data <= "000000000000";
      when "001111010001110" => color_data <= "000000000000";
      when "001111010001111" => color_data <= "000000000000";
      when "001111010010000" => color_data <= "000000000000";
      when "001111010010001" => color_data <= "000000000000";
      when "001111010010010" => color_data <= "110010010000";
      when "001111010010011" => color_data <= "111111000000";
      when "001111010010100" => color_data <= "111111000000";
      when "001111010010101" => color_data <= "110010010001";
      when "001111010010110" => color_data <= "000000000000";
      when "001111010010111" => color_data <= "000000000000";
      when "001111010011000" => color_data <= "000000000000";
      when "001111010011001" => color_data <= "000000000000";
      when "001111010011010" => color_data <= "000000000000";
      when "001111010011011" => color_data <= "000000000000";
      when "001111010011100" => color_data <= "000000000000";
      when "001111010011101" => color_data <= "001100110010";
      when "001111010011110" => color_data <= "110110110000";
      when "001111010011111" => color_data <= "111111010001";
      when "001111010100000" => color_data <= "111111101000";
      when "001111010100001" => color_data <= "111111010011";
      when "001111010100010" => color_data <= "111111010000";
      when "001111010100011" => color_data <= "111111010000";
      when "001111010100100" => color_data <= "111111010000";
      when "001111010100101" => color_data <= "111111010011";
      when "001111010100110" => color_data <= "111111101000";
      when "001111010100111" => color_data <= "111111100111";
      when "001111010101000" => color_data <= "111111100111";
      when "001111010101001" => color_data <= "111111100111";
      when "001111010101010" => color_data <= "111111100111";
      when "001111010101011" => color_data <= "111111100111";
      when "001111010101100" => color_data <= "111111100111";
      when "001111010101101" => color_data <= "111111100111";
      when "001111010101110" => color_data <= "111111100111";
      when "001111010101111" => color_data <= "111111100111";
      when "001111010110000" => color_data <= "111111100111";
      when "001111010110001" => color_data <= "111111100111";
      when "001111010110010" => color_data <= "111111100111";
      when "001111010110011" => color_data <= "111111100111";
      when "001111010110100" => color_data <= "111111100111";
      when "001111010110101" => color_data <= "111111100111";
      when "001111010110110" => color_data <= "111111100111";
      when "001111010110111" => color_data <= "111111100111";
      when "001111010111000" => color_data <= "111111100111";
      when "001111010111001" => color_data <= "111111100111";
      when "001111010111010" => color_data <= "111111100111";
      when "001111010111011" => color_data <= "111111100111";
      when "001111010111100" => color_data <= "111111100110";
      when "001111010111101" => color_data <= "111111101000";
      when "001111010111110" => color_data <= "111111100101";
      when "001111010111111" => color_data <= "111111010000";
      when "001111011000000" => color_data <= "111111000000";
      when "001111011000001" => color_data <= "111111010000";
      when "001111011000010" => color_data <= "111111010000";
      when "001111011000011" => color_data <= "111111010001";
      when "001111011000100" => color_data <= "111111010000";
      when "001111011000101" => color_data <= "110010100000";
      when "001111011000110" => color_data <= "011001100011";
      when "001111011000111" => color_data <= "000000000000";
      when "001111011001000" => color_data <= "000000000000";
      when "001111011001001" => color_data <= "000000000000";
      when "001111011001010" => color_data <= "000000000000";
      when "001111011001011" => color_data <= "000000000000";
      when "001111011001100" => color_data <= "000000000000";
      when "001111011001101" => color_data <= "000000000000";
      when "001111011001110" => color_data <= "000000000000";
      when "001111011001111" => color_data <= "000000000000";
      when "001111011010000" => color_data <= "000000000000";
      when "001111011010001" => color_data <= "010000110010";
      when "001111011010010" => color_data <= "110110100000";
      when "001111011010011" => color_data <= "111111000001";
      when "001111011010100" => color_data <= "110110100000";
      when "001111011010101" => color_data <= "011101100011";
      when "001111011010110" => color_data <= "000000000000";
      when "001111011010111" => color_data <= "000000000000";
      when "001111011011000" => color_data <= "000000000000";
      when "001111011011001" => color_data <= "000000000000";
      when "001111011011010" => color_data <= "000000000000";
      when "001111011011011" => color_data <= "000000000000";
      when "001111011011100" => color_data <= "000000000000";
      when "001111011011101" => color_data <= "000000000000";
      when "001111011011110" => color_data <= "000000000000";
      when "001111011011111" => color_data <= "000000000000";
      when "001111011100000" => color_data <= "000000000000";
      when "001111011100001" => color_data <= "000000000000";
      when "001111011100010" => color_data <= "000000000000";
      when "001111011100011" => color_data <= "000000000000";
      when "001111100000000" => color_data <= "000000000000";
      when "001111100000001" => color_data <= "000000000000";
      when "001111100000010" => color_data <= "000000000000";
      when "001111100000011" => color_data <= "000000000000";
      when "001111100000100" => color_data <= "000000000000";
      when "001111100000101" => color_data <= "000000000000";
      when "001111100000110" => color_data <= "000000000000";
      when "001111100000111" => color_data <= "000000000000";
      when "001111100001000" => color_data <= "000000000000";
      when "001111100001001" => color_data <= "000000000000";
      when "001111100001010" => color_data <= "000000000000";
      when "001111100001011" => color_data <= "000000000000";
      when "001111100001100" => color_data <= "000000000000";
      when "001111100001101" => color_data <= "000000000000";
      when "001111100001110" => color_data <= "000000000000";
      when "001111100001111" => color_data <= "000000000000";
      when "001111100010000" => color_data <= "000000000000";
      when "001111100010001" => color_data <= "000000000000";
      when "001111100010010" => color_data <= "010001000010";
      when "001111100010011" => color_data <= "110110100000";
      when "001111100010100" => color_data <= "111111000001";
      when "001111100010101" => color_data <= "110110100000";
      when "001111100010110" => color_data <= "011101100011";
      when "001111100010111" => color_data <= "000000000000";
      when "001111100011000" => color_data <= "000000000000";
      when "001111100011001" => color_data <= "000000000000";
      when "001111100011010" => color_data <= "000000000000";
      when "001111100011011" => color_data <= "000000000000";
      when "001111100011100" => color_data <= "000000000000";
      when "001111100011101" => color_data <= "000000000000";
      when "001111100011110" => color_data <= "001000100001";
      when "001111100011111" => color_data <= "110110110000";
      when "001111100100000" => color_data <= "111111000000";
      when "001111100100001" => color_data <= "111111010000";
      when "001111100100010" => color_data <= "111111010000";
      when "001111100100011" => color_data <= "111111010001";
      when "001111100100100" => color_data <= "111111010000";
      when "001111100100101" => color_data <= "111111010000";
      when "001111100100110" => color_data <= "111111010100";
      when "001111100100111" => color_data <= "111111101000";
      when "001111100101000" => color_data <= "111111100111";
      when "001111100101001" => color_data <= "111111100111";
      when "001111100101010" => color_data <= "111111100111";
      when "001111100101011" => color_data <= "111111100111";
      when "001111100101100" => color_data <= "111111100111";
      when "001111100101101" => color_data <= "111111100111";
      when "001111100101110" => color_data <= "111111100111";
      when "001111100101111" => color_data <= "111111100111";
      when "001111100110000" => color_data <= "111111100111";
      when "001111100110001" => color_data <= "111111100111";
      when "001111100110010" => color_data <= "111111100111";
      when "001111100110011" => color_data <= "111111100111";
      when "001111100110100" => color_data <= "111111100111";
      when "001111100110101" => color_data <= "111111100111";
      when "001111100110110" => color_data <= "111111100111";
      when "001111100110111" => color_data <= "111111100111";
      when "001111100111000" => color_data <= "111111100111";
      when "001111100111001" => color_data <= "111111100111";
      when "001111100111010" => color_data <= "111111100111";
      when "001111100111011" => color_data <= "111111100111";
      when "001111100111100" => color_data <= "111111100111";
      when "001111100111101" => color_data <= "111111100111";
      when "001111100111110" => color_data <= "111111010001";
      when "001111100111111" => color_data <= "111111010000";
      when "001111101000000" => color_data <= "111111010000";
      when "001111101000001" => color_data <= "111111010000";
      when "001111101000010" => color_data <= "111111010000";
      when "001111101000011" => color_data <= "111111010000";
      when "001111101000100" => color_data <= "110110110000";
      when "001111101000101" => color_data <= "101110010001";
      when "001111101000110" => color_data <= "000000000000";
      when "001111101000111" => color_data <= "000000000000";
      when "001111101001000" => color_data <= "000000000000";
      when "001111101001001" => color_data <= "000000000000";
      when "001111101001010" => color_data <= "000000000000";
      when "001111101001011" => color_data <= "000000000000";
      when "001111101001100" => color_data <= "000000000000";
      when "001111101001101" => color_data <= "000000000000";
      when "001111101001110" => color_data <= "000000000000";
      when "001111101001111" => color_data <= "000000000000";
      when "001111101010000" => color_data <= "000000000000";
      when "001111101010001" => color_data <= "110010010000";
      when "001111101010010" => color_data <= "111111000000";
      when "001111101010011" => color_data <= "111111000000";
      when "001111101010100" => color_data <= "110010010000";
      when "001111101010101" => color_data <= "000000000000";
      when "001111101010110" => color_data <= "000000000000";
      when "001111101010111" => color_data <= "000000000000";
      when "001111101011000" => color_data <= "000000000000";
      when "001111101011001" => color_data <= "000000000000";
      when "001111101011010" => color_data <= "000000000000";
      when "001111101011011" => color_data <= "000000000000";
      when "001111101011100" => color_data <= "000000000000";
      when "001111101011101" => color_data <= "000000000000";
      when "001111101011110" => color_data <= "000000000000";
      when "001111101011111" => color_data <= "000000000000";
      when "001111101100000" => color_data <= "000000000000";
      when "001111101100001" => color_data <= "000000000000";
      when "001111101100010" => color_data <= "000000000000";
      when "001111101100011" => color_data <= "000000000000";
      when "001111110000000" => color_data <= "000000000000";
      when "001111110000001" => color_data <= "000000000000";
      when "001111110000010" => color_data <= "000000000000";
      when "001111110000011" => color_data <= "000000000000";
      when "001111110000100" => color_data <= "000000000000";
      when "001111110000101" => color_data <= "000000000000";
      when "001111110000110" => color_data <= "000000000000";
      when "001111110000111" => color_data <= "000000000000";
      when "001111110001000" => color_data <= "000000000000";
      when "001111110001001" => color_data <= "000000000000";
      when "001111110001010" => color_data <= "000000000000";
      when "001111110001011" => color_data <= "000000000000";
      when "001111110001100" => color_data <= "000000000000";
      when "001111110001101" => color_data <= "000000000000";
      when "001111110001110" => color_data <= "000000000000";
      when "001111110001111" => color_data <= "000000000000";
      when "001111110010000" => color_data <= "000000000000";
      when "001111110010001" => color_data <= "000000000000";
      when "001111110010010" => color_data <= "000000000000";
      when "001111110010011" => color_data <= "101010000010";
      when "001111110010100" => color_data <= "111110110000";
      when "001111110010101" => color_data <= "111111000001";
      when "001111110010110" => color_data <= "110110100000";
      when "001111110010111" => color_data <= "000100010001";
      when "001111110011000" => color_data <= "000000000000";
      when "001111110011001" => color_data <= "000000000000";
      when "001111110011010" => color_data <= "000000000000";
      when "001111110011011" => color_data <= "000000000000";
      when "001111110011100" => color_data <= "000000000000";
      when "001111110011101" => color_data <= "000000000000";
      when "001111110011110" => color_data <= "000000000000";
      when "001111110011111" => color_data <= "000000000000";
      when "001111110100000" => color_data <= "101110010001";
      when "001111110100001" => color_data <= "110110110000";
      when "001111110100010" => color_data <= "111111010000";
      when "001111110100011" => color_data <= "111111010001";
      when "001111110100100" => color_data <= "111111010000";
      when "001111110100101" => color_data <= "111111010000";
      when "001111110100110" => color_data <= "111111010000";
      when "001111110100111" => color_data <= "111111100110";
      when "001111110101000" => color_data <= "111111101000";
      when "001111110101001" => color_data <= "111111100110";
      when "001111110101010" => color_data <= "111111100111";
      when "001111110101011" => color_data <= "111111100111";
      when "001111110101100" => color_data <= "111111100111";
      when "001111110101101" => color_data <= "111111100111";
      when "001111110101110" => color_data <= "111111100111";
      when "001111110101111" => color_data <= "111111100111";
      when "001111110110000" => color_data <= "111111100111";
      when "001111110110001" => color_data <= "111111100111";
      when "001111110110010" => color_data <= "111111100111";
      when "001111110110011" => color_data <= "111111100111";
      when "001111110110100" => color_data <= "111111100111";
      when "001111110110101" => color_data <= "111111100111";
      when "001111110110110" => color_data <= "111111100111";
      when "001111110110111" => color_data <= "111111100111";
      when "001111110111000" => color_data <= "111111100111";
      when "001111110111001" => color_data <= "111111100111";
      when "001111110111010" => color_data <= "111111100111";
      when "001111110111011" => color_data <= "111111100111";
      when "001111110111100" => color_data <= "111111101000";
      when "001111110111101" => color_data <= "111111010011";
      when "001111110111110" => color_data <= "111111010000";
      when "001111110111111" => color_data <= "111111010000";
      when "001111111000000" => color_data <= "111111010000";
      when "001111111000001" => color_data <= "111111010000";
      when "001111111000010" => color_data <= "111111010000";
      when "001111111000011" => color_data <= "110110110000";
      when "001111111000100" => color_data <= "100001110010";
      when "001111111000101" => color_data <= "000000000000";
      when "001111111000110" => color_data <= "000000000000";
      when "001111111000111" => color_data <= "000000000000";
      when "001111111001000" => color_data <= "000000000000";
      when "001111111001001" => color_data <= "000000000000";
      when "001111111001010" => color_data <= "000000000000";
      when "001111111001011" => color_data <= "000000000000";
      when "001111111001100" => color_data <= "000000000000";
      when "001111111001101" => color_data <= "000000000000";
      when "001111111001110" => color_data <= "000000000000";
      when "001111111001111" => color_data <= "000000000000";
      when "001111111010000" => color_data <= "100001110010";
      when "001111111010001" => color_data <= "110110100000";
      when "001111111010010" => color_data <= "111111000001";
      when "001111111010011" => color_data <= "110110100000";
      when "001111111010100" => color_data <= "001100110010";
      when "001111111010101" => color_data <= "000000000000";
      when "001111111010110" => color_data <= "000000000000";
      when "001111111010111" => color_data <= "000000000000";
      when "001111111011000" => color_data <= "000000000000";
      when "001111111011001" => color_data <= "000000000000";
      when "001111111011010" => color_data <= "000000000000";
      when "001111111011011" => color_data <= "000000000000";
      when "001111111011100" => color_data <= "000000000000";
      when "001111111011101" => color_data <= "000000000000";
      when "001111111011110" => color_data <= "000000000000";
      when "001111111011111" => color_data <= "000000000000";
      when "001111111100000" => color_data <= "000000000000";
      when "001111111100001" => color_data <= "000000000000";
      when "001111111100010" => color_data <= "000000000000";
      when "001111111100011" => color_data <= "000000000000";
      when "010000000000000" => color_data <= "000000000000";
      when "010000000000001" => color_data <= "000000000000";
      when "010000000000010" => color_data <= "000000000000";
      when "010000000000011" => color_data <= "000000000000";
      when "010000000000100" => color_data <= "000000000000";
      when "010000000000101" => color_data <= "000000000000";
      when "010000000000110" => color_data <= "000000000000";
      when "010000000000111" => color_data <= "000000000000";
      when "010000000001000" => color_data <= "000000000000";
      when "010000000001001" => color_data <= "000000000000";
      when "010000000001010" => color_data <= "000000000000";
      when "010000000001011" => color_data <= "000000000000";
      when "010000000001100" => color_data <= "000000000000";
      when "010000000001101" => color_data <= "000000000000";
      when "010000000001110" => color_data <= "000000000000";
      when "010000000001111" => color_data <= "000000000000";
      when "010000000010000" => color_data <= "000000000000";
      when "010000000010001" => color_data <= "000000000000";
      when "010000000010010" => color_data <= "000000000000";
      when "010000000010011" => color_data <= "000000000000";
      when "010000000010100" => color_data <= "110110100000";
      when "010000000010101" => color_data <= "111111000000";
      when "010000000010110" => color_data <= "111110110000";
      when "010000000010111" => color_data <= "101110010001";
      when "010000000011000" => color_data <= "000000000000";
      when "010000000011001" => color_data <= "000000000000";
      when "010000000011010" => color_data <= "000000000000";
      when "010000000011011" => color_data <= "000000000000";
      when "010000000011100" => color_data <= "000000000000";
      when "010000000011101" => color_data <= "000000000000";
      when "010000000011110" => color_data <= "000000000000";
      when "010000000011111" => color_data <= "000000000000";
      when "010000000100000" => color_data <= "000000000000";
      when "010000000100001" => color_data <= "011001010011";
      when "010000000100010" => color_data <= "110110110000";
      when "010000000100011" => color_data <= "111111000000";
      when "010000000100100" => color_data <= "111111010000";
      when "010000000100101" => color_data <= "111111010001";
      when "010000000100110" => color_data <= "111111010000";
      when "010000000100111" => color_data <= "111111010001";
      when "010000000101000" => color_data <= "111111100111";
      when "010000000101001" => color_data <= "111111100111";
      when "010000000101010" => color_data <= "111111100110";
      when "010000000101011" => color_data <= "111111100111";
      when "010000000101100" => color_data <= "111111100111";
      when "010000000101101" => color_data <= "111111100111";
      when "010000000101110" => color_data <= "111111100111";
      when "010000000101111" => color_data <= "111111100111";
      when "010000000110000" => color_data <= "111111100111";
      when "010000000110001" => color_data <= "111111100111";
      when "010000000110010" => color_data <= "111111100111";
      when "010000000110011" => color_data <= "111111100111";
      when "010000000110100" => color_data <= "111111100111";
      when "010000000110101" => color_data <= "111111100111";
      when "010000000110110" => color_data <= "111111100111";
      when "010000000110111" => color_data <= "111111100111";
      when "010000000111000" => color_data <= "111111100111";
      when "010000000111001" => color_data <= "111111100111";
      when "010000000111010" => color_data <= "111111100110";
      when "010000000111011" => color_data <= "111111101000";
      when "010000000111100" => color_data <= "111111100101";
      when "010000000111101" => color_data <= "111111010000";
      when "010000000111110" => color_data <= "111111010000";
      when "010000000111111" => color_data <= "111111010001";
      when "010000001000000" => color_data <= "111111010000";
      when "010000001000001" => color_data <= "110110110000";
      when "010000001000010" => color_data <= "110010100000";
      when "010000001000011" => color_data <= "010000110010";
      when "010000001000100" => color_data <= "000000000000";
      when "010000001000101" => color_data <= "000000000000";
      when "010000001000110" => color_data <= "000000000000";
      when "010000001000111" => color_data <= "000000000000";
      when "010000001001000" => color_data <= "000000000000";
      when "010000001001001" => color_data <= "000000000000";
      when "010000001001010" => color_data <= "000000000000";
      when "010000001001011" => color_data <= "000000000000";
      when "010000001001100" => color_data <= "000000000000";
      when "010000001001101" => color_data <= "000000000000";
      when "010000001001110" => color_data <= "000000000000";
      when "010000001001111" => color_data <= "001100100010";
      when "010000001010000" => color_data <= "110110100000";
      when "010000001010001" => color_data <= "111111000001";
      when "010000001010010" => color_data <= "110110100000";
      when "010000001010011" => color_data <= "100110000010";
      when "010000001010100" => color_data <= "000000000000";
      when "010000001010101" => color_data <= "000000000000";
      when "010000001010110" => color_data <= "000000000000";
      when "010000001010111" => color_data <= "000000000000";
      when "010000001011000" => color_data <= "000000000000";
      when "010000001011001" => color_data <= "000000000000";
      when "010000001011010" => color_data <= "000000000000";
      when "010000001011011" => color_data <= "000000000000";
      when "010000001011100" => color_data <= "000000000000";
      when "010000001011101" => color_data <= "000000000000";
      when "010000001011110" => color_data <= "000000000000";
      when "010000001011111" => color_data <= "000000000000";
      when "010000001100000" => color_data <= "000000000000";
      when "010000001100001" => color_data <= "000000000000";
      when "010000001100010" => color_data <= "000000000000";
      when "010000001100011" => color_data <= "000000000000";
      when "010000010000000" => color_data <= "000000000000";
      when "010000010000001" => color_data <= "000000000000";
      when "010000010000010" => color_data <= "000000000000";
      when "010000010000011" => color_data <= "000000000000";
      when "010000010000100" => color_data <= "000000000000";
      when "010000010000101" => color_data <= "000000000000";
      when "010000010000110" => color_data <= "000000000000";
      when "010000010000111" => color_data <= "000000000000";
      when "010000010001000" => color_data <= "000000000000";
      when "010000010001001" => color_data <= "000000000000";
      when "010000010001010" => color_data <= "000000000000";
      when "010000010001011" => color_data <= "000000000000";
      when "010000010001100" => color_data <= "000000000000";
      when "010000010001101" => color_data <= "000000000000";
      when "010000010001110" => color_data <= "000000000000";
      when "010000010001111" => color_data <= "000000000000";
      when "010000010010000" => color_data <= "000000000000";
      when "010000010010001" => color_data <= "000000000000";
      when "010000010010010" => color_data <= "000000000000";
      when "010000010010011" => color_data <= "000000000000";
      when "010000010010100" => color_data <= "010101010011";
      when "010000010010101" => color_data <= "110110100000";
      when "010000010010110" => color_data <= "111111000001";
      when "010000010010111" => color_data <= "110110100000";
      when "010000010011000" => color_data <= "011101100011";
      when "010000010011001" => color_data <= "000000000000";
      when "010000010011010" => color_data <= "000000000000";
      when "010000010011011" => color_data <= "000000000000";
      when "010000010011100" => color_data <= "000000000000";
      when "010000010011101" => color_data <= "000000000000";
      when "010000010011110" => color_data <= "000000000000";
      when "010000010011111" => color_data <= "000000000000";
      when "010000010100000" => color_data <= "000000000000";
      when "010000010100001" => color_data <= "000000000000";
      when "010000010100010" => color_data <= "000100010001";
      when "010000010100011" => color_data <= "101010000010";
      when "010000010100100" => color_data <= "110110110000";
      when "010000010100101" => color_data <= "111111000000";
      when "010000010100110" => color_data <= "111111010000";
      when "010000010100111" => color_data <= "111111010000";
      when "010000010101000" => color_data <= "111111010010";
      when "010000010101001" => color_data <= "111111101000";
      when "010000010101010" => color_data <= "111111100111";
      when "010000010101011" => color_data <= "111111100111";
      when "010000010101100" => color_data <= "111111100111";
      when "010000010101101" => color_data <= "111111100111";
      when "010000010101110" => color_data <= "111111100111";
      when "010000010101111" => color_data <= "111111100111";
      when "010000010110000" => color_data <= "111111100111";
      when "010000010110001" => color_data <= "111111100111";
      when "010000010110010" => color_data <= "111111100111";
      when "010000010110011" => color_data <= "111111100111";
      when "010000010110100" => color_data <= "111111100111";
      when "010000010110101" => color_data <= "111111100111";
      when "010000010110110" => color_data <= "111111100111";
      when "010000010110111" => color_data <= "111111100111";
      when "010000010111000" => color_data <= "111111100111";
      when "010000010111001" => color_data <= "111111100110";
      when "010000010111010" => color_data <= "111111100111";
      when "010000010111011" => color_data <= "111111100111";
      when "010000010111100" => color_data <= "111111010000";
      when "010000010111101" => color_data <= "111111010000";
      when "010000010111110" => color_data <= "111111010000";
      when "010000010111111" => color_data <= "111111000000";
      when "010000011000000" => color_data <= "110110110000";
      when "010000011000001" => color_data <= "100001110010";
      when "010000011000010" => color_data <= "000000000000";
      when "010000011000011" => color_data <= "000000000000";
      when "010000011000100" => color_data <= "000000000000";
      when "010000011000101" => color_data <= "000000000000";
      when "010000011000110" => color_data <= "000000000000";
      when "010000011000111" => color_data <= "000000000000";
      when "010000011001000" => color_data <= "000000000000";
      when "010000011001001" => color_data <= "000000000000";
      when "010000011001010" => color_data <= "000000000000";
      when "010000011001011" => color_data <= "000000000000";
      when "010000011001100" => color_data <= "000000000000";
      when "010000011001101" => color_data <= "000000000000";
      when "010000011001110" => color_data <= "000000000000";
      when "010000011001111" => color_data <= "110010010000";
      when "010000011010000" => color_data <= "111111000000";
      when "010000011010001" => color_data <= "111111000000";
      when "010000011010010" => color_data <= "110110100000";
      when "010000011010011" => color_data <= "000000000000";
      when "010000011010100" => color_data <= "000000000000";
      when "010000011010101" => color_data <= "000000000000";
      when "010000011010110" => color_data <= "000000000000";
      when "010000011010111" => color_data <= "000000000000";
      when "010000011011000" => color_data <= "000000000000";
      when "010000011011001" => color_data <= "000000000000";
      when "010000011011010" => color_data <= "000000000000";
      when "010000011011011" => color_data <= "000000000000";
      when "010000011011100" => color_data <= "000000000000";
      when "010000011011101" => color_data <= "000000000000";
      when "010000011011110" => color_data <= "000000000000";
      when "010000011011111" => color_data <= "000000000000";
      when "010000011100000" => color_data <= "000000000000";
      when "010000011100001" => color_data <= "000000000000";
      when "010000011100010" => color_data <= "000000000000";
      when "010000011100011" => color_data <= "000000000000";
      when "010000100000000" => color_data <= "000000000000";
      when "010000100000001" => color_data <= "000000000000";
      when "010000100000010" => color_data <= "000000000000";
      when "010000100000011" => color_data <= "000000000000";
      when "010000100000100" => color_data <= "000000000000";
      when "010000100000101" => color_data <= "000000000000";
      when "010000100000110" => color_data <= "000000000000";
      when "010000100000111" => color_data <= "000000000000";
      when "010000100001000" => color_data <= "000000000000";
      when "010000100001001" => color_data <= "000000000000";
      when "010000100001010" => color_data <= "000000000000";
      when "010000100001011" => color_data <= "000000000000";
      when "010000100001100" => color_data <= "000000000000";
      when "010000100001101" => color_data <= "000000000000";
      when "010000100001110" => color_data <= "000000000000";
      when "010000100001111" => color_data <= "000000000000";
      when "010000100010000" => color_data <= "000000000000";
      when "010000100010001" => color_data <= "000000000000";
      when "010000100010010" => color_data <= "000000000000";
      when "010000100010011" => color_data <= "000000000000";
      when "010000100010100" => color_data <= "000000000000";
      when "010000100010101" => color_data <= "100110000010";
      when "010000100010110" => color_data <= "111110110000";
      when "010000100010111" => color_data <= "111111000001";
      when "010000100011000" => color_data <= "110110100000";
      when "010000100011001" => color_data <= "001100110010";
      when "010000100011010" => color_data <= "000000000000";
      when "010000100011011" => color_data <= "000000000000";
      when "010000100011100" => color_data <= "000000000000";
      when "010000100011101" => color_data <= "000000000000";
      when "010000100011110" => color_data <= "000000000000";
      when "010000100011111" => color_data <= "000000000000";
      when "010000100100000" => color_data <= "000000000000";
      when "010000100100001" => color_data <= "000000000000";
      when "010000100100010" => color_data <= "000000000000";
      when "010000100100011" => color_data <= "000000000000";
      when "010000100100100" => color_data <= "001100110010";
      when "010000100100101" => color_data <= "101010000010";
      when "010000100100110" => color_data <= "110110110000";
      when "010000100100111" => color_data <= "111111000000";
      when "010000100101000" => color_data <= "111111000000";
      when "010000100101001" => color_data <= "111111010100";
      when "010000100101010" => color_data <= "111111101000";
      when "010000100101011" => color_data <= "111111100111";
      when "010000100101100" => color_data <= "111111100111";
      when "010000100101101" => color_data <= "111111100111";
      when "010000100101110" => color_data <= "111111100111";
      when "010000100101111" => color_data <= "111111100111";
      when "010000100110000" => color_data <= "111111100111";
      when "010000100110001" => color_data <= "111111100111";
      when "010000100110010" => color_data <= "111111100111";
      when "010000100110011" => color_data <= "111111100111";
      when "010000100110100" => color_data <= "111111100111";
      when "010000100110101" => color_data <= "111111100111";
      when "010000100110110" => color_data <= "111111100111";
      when "010000100110111" => color_data <= "111111100111";
      when "010000100111000" => color_data <= "111111100110";
      when "010000100111001" => color_data <= "111111100111";
      when "010000100111010" => color_data <= "111111101000";
      when "010000100111011" => color_data <= "111111010001";
      when "010000100111100" => color_data <= "111111000000";
      when "010000100111101" => color_data <= "111111000000";
      when "010000100111110" => color_data <= "110110110000";
      when "010000100111111" => color_data <= "100001110010";
      when "010000101000000" => color_data <= "000100010001";
      when "010000101000001" => color_data <= "000000000000";
      when "010000101000010" => color_data <= "000000000000";
      when "010000101000011" => color_data <= "000000000000";
      when "010000101000100" => color_data <= "000000000000";
      when "010000101000101" => color_data <= "000000000000";
      when "010000101000110" => color_data <= "000000000000";
      when "010000101000111" => color_data <= "000000000000";
      when "010000101001000" => color_data <= "000000000000";
      when "010000101001001" => color_data <= "000000000000";
      when "010000101001010" => color_data <= "000000000000";
      when "010000101001011" => color_data <= "000000000000";
      when "010000101001100" => color_data <= "000000000000";
      when "010000101001101" => color_data <= "000000000000";
      when "010000101001110" => color_data <= "100110000010";
      when "010000101001111" => color_data <= "110110100000";
      when "010000101010000" => color_data <= "111111000000";
      when "010000101010001" => color_data <= "110110100000";
      when "010000101010010" => color_data <= "001000100010";
      when "010000101010011" => color_data <= "000000000000";
      when "010000101010100" => color_data <= "000000000000";
      when "010000101010101" => color_data <= "000000000000";
      when "010000101010110" => color_data <= "000000000000";
      when "010000101010111" => color_data <= "000000000000";
      when "010000101011000" => color_data <= "000000000000";
      when "010000101011001" => color_data <= "000000000000";
      when "010000101011010" => color_data <= "000000000000";
      when "010000101011011" => color_data <= "000000000000";
      when "010000101011100" => color_data <= "000000000000";
      when "010000101011101" => color_data <= "000000000000";
      when "010000101011110" => color_data <= "000000000000";
      when "010000101011111" => color_data <= "000000000000";
      when "010000101100000" => color_data <= "000000000000";
      when "010000101100001" => color_data <= "000000000000";
      when "010000101100010" => color_data <= "000000000000";
      when "010000101100011" => color_data <= "000000000000";
      when "010000110000000" => color_data <= "000000000000";
      when "010000110000001" => color_data <= "000000000000";
      when "010000110000010" => color_data <= "000000000000";
      when "010000110000011" => color_data <= "000000000000";
      when "010000110000100" => color_data <= "000000000000";
      when "010000110000101" => color_data <= "000000000000";
      when "010000110000110" => color_data <= "000000000000";
      when "010000110000111" => color_data <= "000000000000";
      when "010000110001000" => color_data <= "000000000000";
      when "010000110001001" => color_data <= "000000000000";
      when "010000110001010" => color_data <= "000000000000";
      when "010000110001011" => color_data <= "000000000000";
      when "010000110001100" => color_data <= "000000000000";
      when "010000110001101" => color_data <= "000000000000";
      when "010000110001110" => color_data <= "000000000000";
      when "010000110001111" => color_data <= "000000000000";
      when "010000110010000" => color_data <= "000000000000";
      when "010000110010001" => color_data <= "000000000000";
      when "010000110010010" => color_data <= "000000000000";
      when "010000110010011" => color_data <= "000000000000";
      when "010000110010100" => color_data <= "000000000000";
      when "010000110010101" => color_data <= "000000000000";
      when "010000110010110" => color_data <= "110110100000";
      when "010000110010111" => color_data <= "111111000000";
      when "010000110011000" => color_data <= "111111000000";
      when "010000110011001" => color_data <= "110010100000";
      when "010000110011010" => color_data <= "000000000000";
      when "010000110011011" => color_data <= "000000000000";
      when "010000110011100" => color_data <= "000000000000";
      when "010000110011101" => color_data <= "000000000000";
      when "010000110011110" => color_data <= "000000000000";
      when "010000110011111" => color_data <= "000000000000";
      when "010000110100000" => color_data <= "000000000000";
      when "010000110100001" => color_data <= "000000000000";
      when "010000110100010" => color_data <= "000000000000";
      when "010000110100011" => color_data <= "000000000000";
      when "010000110100100" => color_data <= "000000000000";
      when "010000110100101" => color_data <= "000000000000";
      when "010000110100110" => color_data <= "001000100001";
      when "010000110100111" => color_data <= "100001110010";
      when "010000110101000" => color_data <= "110110100000";
      when "010000110101001" => color_data <= "110110110000";
      when "010000110101010" => color_data <= "111111010011";
      when "010000110101011" => color_data <= "111111100111";
      when "010000110101100" => color_data <= "111111100111";
      when "010000110101101" => color_data <= "111111100111";
      when "010000110101110" => color_data <= "111111100111";
      when "010000110101111" => color_data <= "111111100111";
      when "010000110110000" => color_data <= "111111100111";
      when "010000110110001" => color_data <= "111111100111";
      when "010000110110010" => color_data <= "111111100111";
      when "010000110110011" => color_data <= "111111100111";
      when "010000110110100" => color_data <= "111111100111";
      when "010000110110101" => color_data <= "111111100111";
      when "010000110110110" => color_data <= "111111100111";
      when "010000110110111" => color_data <= "111111100111";
      when "010000110111000" => color_data <= "111111100111";
      when "010000110111001" => color_data <= "111111100110";
      when "010000110111010" => color_data <= "111111010000";
      when "010000110111011" => color_data <= "110110110000";
      when "010000110111100" => color_data <= "101110100001";
      when "010000110111101" => color_data <= "011101100011";
      when "010000110111110" => color_data <= "000000000000";
      when "010000110111111" => color_data <= "000000000000";
      when "010000111000000" => color_data <= "000000000000";
      when "010000111000001" => color_data <= "000000000000";
      when "010000111000010" => color_data <= "000000000000";
      when "010000111000011" => color_data <= "000000000000";
      when "010000111000100" => color_data <= "000000000000";
      when "010000111000101" => color_data <= "000000000000";
      when "010000111000110" => color_data <= "000000000000";
      when "010000111000111" => color_data <= "000000000000";
      when "010000111001000" => color_data <= "000000000000";
      when "010000111001001" => color_data <= "000000000000";
      when "010000111001010" => color_data <= "000000000000";
      when "010000111001011" => color_data <= "000000000000";
      when "010000111001100" => color_data <= "000000000000";
      when "010000111001101" => color_data <= "011001010011";
      when "010000111001110" => color_data <= "110110100000";
      when "010000111001111" => color_data <= "111111000001";
      when "010000111010000" => color_data <= "110110100000";
      when "010000111010001" => color_data <= "011101100011";
      when "010000111010010" => color_data <= "000000000000";
      when "010000111010011" => color_data <= "000000000000";
      when "010000111010100" => color_data <= "000000000000";
      when "010000111010101" => color_data <= "000000000000";
      when "010000111010110" => color_data <= "000000000000";
      when "010000111010111" => color_data <= "000000000000";
      when "010000111011000" => color_data <= "000000000000";
      when "010000111011001" => color_data <= "000000000000";
      when "010000111011010" => color_data <= "000000000000";
      when "010000111011011" => color_data <= "000000000000";
      when "010000111011100" => color_data <= "000000000000";
      when "010000111011101" => color_data <= "000000000000";
      when "010000111011110" => color_data <= "000000000000";
      when "010000111011111" => color_data <= "000000000000";
      when "010000111100000" => color_data <= "000000000000";
      when "010000111100001" => color_data <= "000000000000";
      when "010000111100010" => color_data <= "000000000000";
      when "010000111100011" => color_data <= "000000000000";
      when "010001000000000" => color_data <= "000000000000";
      when "010001000000001" => color_data <= "000000000000";
      when "010001000000010" => color_data <= "000000000000";
      when "010001000000011" => color_data <= "000000000000";
      when "010001000000100" => color_data <= "000000000000";
      when "010001000000101" => color_data <= "000000000000";
      when "010001000000110" => color_data <= "000000000000";
      when "010001000000111" => color_data <= "000000000000";
      when "010001000001000" => color_data <= "000000000000";
      when "010001000001001" => color_data <= "000000000000";
      when "010001000001010" => color_data <= "000000000000";
      when "010001000001011" => color_data <= "000000000000";
      when "010001000001100" => color_data <= "000000000000";
      when "010001000001101" => color_data <= "000000000000";
      when "010001000001110" => color_data <= "000000000000";
      when "010001000001111" => color_data <= "000000000000";
      when "010001000010000" => color_data <= "000000000000";
      when "010001000010001" => color_data <= "000000000000";
      when "010001000010010" => color_data <= "000000000000";
      when "010001000010011" => color_data <= "000000000000";
      when "010001000010100" => color_data <= "000000000000";
      when "010001000010101" => color_data <= "000000000000";
      when "010001000010110" => color_data <= "001000100010";
      when "010001000010111" => color_data <= "110110100000";
      when "010001000011000" => color_data <= "111111000000";
      when "010001000011001" => color_data <= "110110100000";
      when "010001000011010" => color_data <= "101010000001";
      when "010001000011011" => color_data <= "000000000000";
      when "010001000011100" => color_data <= "000000000000";
      when "010001000011101" => color_data <= "000000000000";
      when "010001000011110" => color_data <= "000000000000";
      when "010001000011111" => color_data <= "000000000000";
      when "010001000100000" => color_data <= "000000000000";
      when "010001000100001" => color_data <= "000000000000";
      when "010001000100010" => color_data <= "000000000000";
      when "010001000100011" => color_data <= "000000000000";
      when "010001000100100" => color_data <= "000000000000";
      when "010001000100101" => color_data <= "000000000000";
      when "010001000100110" => color_data <= "000000000000";
      when "010001000100111" => color_data <= "000000000000";
      when "010001000101000" => color_data <= "000000000000";
      when "010001000101001" => color_data <= "010001000010";
      when "010001000101010" => color_data <= "011001100011";
      when "010001000101011" => color_data <= "011101110011";
      when "010001000101100" => color_data <= "100010000010";
      when "010001000101101" => color_data <= "111111010101";
      when "010001000101110" => color_data <= "111111010100";
      when "010001000101111" => color_data <= "111111010100";
      when "010001000110000" => color_data <= "111111010101";
      when "010001000110001" => color_data <= "111111100101";
      when "010001000110010" => color_data <= "111111100101";
      when "010001000110011" => color_data <= "111111100101";
      when "010001000110100" => color_data <= "111111010101";
      when "010001000110101" => color_data <= "111111010100";
      when "010001000110110" => color_data <= "111111010100";
      when "010001000110111" => color_data <= "111111100101";
      when "010001000111000" => color_data <= "100001110010";
      when "010001000111001" => color_data <= "100001110010";
      when "010001000111010" => color_data <= "011101100011";
      when "010001000111011" => color_data <= "001000100010";
      when "010001000111100" => color_data <= "000000000000";
      when "010001000111101" => color_data <= "000000000000";
      when "010001000111110" => color_data <= "000000000000";
      when "010001000111111" => color_data <= "000000000000";
      when "010001001000000" => color_data <= "000000000000";
      when "010001001000001" => color_data <= "000000000000";
      when "010001001000010" => color_data <= "000000000000";
      when "010001001000011" => color_data <= "000000000000";
      when "010001001000100" => color_data <= "000000000000";
      when "010001001000101" => color_data <= "000000000000";
      when "010001001000110" => color_data <= "000000000000";
      when "010001001000111" => color_data <= "000000000000";
      when "010001001001000" => color_data <= "000000000000";
      when "010001001001001" => color_data <= "000000000000";
      when "010001001001010" => color_data <= "000000000000";
      when "010001001001011" => color_data <= "000000000000";
      when "010001001001100" => color_data <= "001100110010";
      when "010001001001101" => color_data <= "110110100000";
      when "010001001001110" => color_data <= "111111000000";
      when "010001001001111" => color_data <= "110110100000";
      when "010001001010000" => color_data <= "101010000010";
      when "010001001010001" => color_data <= "000000000000";
      when "010001001010010" => color_data <= "000000000000";
      when "010001001010011" => color_data <= "000000000000";
      when "010001001010100" => color_data <= "000000000000";
      when "010001001010101" => color_data <= "000000000000";
      when "010001001010110" => color_data <= "000000000000";
      when "010001001010111" => color_data <= "000000000000";
      when "010001001011000" => color_data <= "000000000000";
      when "010001001011001" => color_data <= "000000000000";
      when "010001001011010" => color_data <= "000000000000";
      when "010001001011011" => color_data <= "000000000000";
      when "010001001011100" => color_data <= "000000000000";
      when "010001001011101" => color_data <= "000000000000";
      when "010001001011110" => color_data <= "000000000000";
      when "010001001011111" => color_data <= "000000000000";
      when "010001001100000" => color_data <= "000000000000";
      when "010001001100001" => color_data <= "000000000000";
      when "010001001100010" => color_data <= "000000000000";
      when "010001001100011" => color_data <= "000000000000";
      when "010001010000000" => color_data <= "000000000000";
      when "010001010000001" => color_data <= "000000000000";
      when "010001010000010" => color_data <= "000000000000";
      when "010001010000011" => color_data <= "000000000000";
      when "010001010000100" => color_data <= "000000000000";
      when "010001010000101" => color_data <= "000000000000";
      when "010001010000110" => color_data <= "000000000000";
      when "010001010000111" => color_data <= "000000000000";
      when "010001010001000" => color_data <= "000000000000";
      when "010001010001001" => color_data <= "000000000000";
      when "010001010001010" => color_data <= "000000000000";
      when "010001010001011" => color_data <= "000000000000";
      when "010001010001100" => color_data <= "000000000000";
      when "010001010001101" => color_data <= "000000000000";
      when "010001010001110" => color_data <= "000000000000";
      when "010001010001111" => color_data <= "000000000000";
      when "010001010010000" => color_data <= "000000000000";
      when "010001010010001" => color_data <= "000000000000";
      when "010001010010010" => color_data <= "000000000000";
      when "010001010010011" => color_data <= "000000000000";
      when "010001010010100" => color_data <= "000000000000";
      when "010001010010101" => color_data <= "000000000000";
      when "010001010010110" => color_data <= "000000000000";
      when "010001010010111" => color_data <= "011001010011";
      when "010001010011000" => color_data <= "110110100000";
      when "010001010011001" => color_data <= "111111000001";
      when "010001010011010" => color_data <= "110110100000";
      when "010001010011011" => color_data <= "100001110010";
      when "010001010011100" => color_data <= "000000000000";
      when "010001010011101" => color_data <= "000000000000";
      when "010001010011110" => color_data <= "000000000000";
      when "010001010011111" => color_data <= "000000000000";
      when "010001010100000" => color_data <= "000000000000";
      when "010001010100001" => color_data <= "000000000000";
      when "010001010100010" => color_data <= "000000000000";
      when "010001010100011" => color_data <= "000000000000";
      when "010001010100100" => color_data <= "000000000000";
      when "010001010100101" => color_data <= "000000000000";
      when "010001010100110" => color_data <= "000000000000";
      when "010001010100111" => color_data <= "000000000000";
      when "010001010101000" => color_data <= "000000000000";
      when "010001010101001" => color_data <= "000000000000";
      when "010001010101010" => color_data <= "000000000000";
      when "010001010101011" => color_data <= "000000000000";
      when "010001010101100" => color_data <= "000100010001";
      when "010001010101101" => color_data <= "000100010001";
      when "010001010101110" => color_data <= "001100110010";
      when "010001010101111" => color_data <= "010001000010";
      when "010001010110000" => color_data <= "011001010011";
      when "010001010110001" => color_data <= "011001010011";
      when "010001010110010" => color_data <= "011001010011";
      when "010001010110011" => color_data <= "011001010011";
      when "010001010110100" => color_data <= "011001010011";
      when "010001010110101" => color_data <= "010001000010";
      when "010001010110110" => color_data <= "001100100010";
      when "010001010110111" => color_data <= "000100010001";
      when "010001010111000" => color_data <= "000100010001";
      when "010001010111001" => color_data <= "000000000000";
      when "010001010111010" => color_data <= "000000000000";
      when "010001010111011" => color_data <= "000000000000";
      when "010001010111100" => color_data <= "000000000000";
      when "010001010111101" => color_data <= "000000000000";
      when "010001010111110" => color_data <= "000000000000";
      when "010001010111111" => color_data <= "000000000000";
      when "010001011000000" => color_data <= "000000000000";
      when "010001011000001" => color_data <= "000000000000";
      when "010001011000010" => color_data <= "000000000000";
      when "010001011000011" => color_data <= "000000000000";
      when "010001011000100" => color_data <= "000000000000";
      when "010001011000101" => color_data <= "000000000000";
      when "010001011000110" => color_data <= "000000000000";
      when "010001011000111" => color_data <= "000000000000";
      when "010001011001000" => color_data <= "000000000000";
      when "010001011001001" => color_data <= "000000000000";
      when "010001011001010" => color_data <= "000000000000";
      when "010001011001011" => color_data <= "000100010001";
      when "010001011001100" => color_data <= "110110100000";
      when "010001011001101" => color_data <= "111111000000";
      when "010001011001110" => color_data <= "111110110000";
      when "010001011001111" => color_data <= "110010100000";
      when "010001011010000" => color_data <= "000000000000";
      when "010001011010001" => color_data <= "000000000000";
      when "010001011010010" => color_data <= "000000000000";
      when "010001011010011" => color_data <= "000000000000";
      when "010001011010100" => color_data <= "000000000000";
      when "010001011010101" => color_data <= "000000000000";
      when "010001011010110" => color_data <= "000000000000";
      when "010001011010111" => color_data <= "000000000000";
      when "010001011011000" => color_data <= "000000000000";
      when "010001011011001" => color_data <= "000000000000";
      when "010001011011010" => color_data <= "000000000000";
      when "010001011011011" => color_data <= "000000000000";
      when "010001011011100" => color_data <= "000000000000";
      when "010001011011101" => color_data <= "000000000000";
      when "010001011011110" => color_data <= "000000000000";
      when "010001011011111" => color_data <= "000000000000";
      when "010001011100000" => color_data <= "000000000000";
      when "010001011100001" => color_data <= "000000000000";
      when "010001011100010" => color_data <= "000000000000";
      when "010001011100011" => color_data <= "000000000000";
      when "010001100000000" => color_data <= "000000000000";
      when "010001100000001" => color_data <= "000000000000";
      when "010001100000010" => color_data <= "000000000000";
      when "010001100000011" => color_data <= "000000000000";
      when "010001100000100" => color_data <= "000000000000";
      when "010001100000101" => color_data <= "000000000000";
      when "010001100000110" => color_data <= "000000000000";
      when "010001100000111" => color_data <= "000000000000";
      when "010001100001000" => color_data <= "000000000000";
      when "010001100001001" => color_data <= "000000000000";
      when "010001100001010" => color_data <= "000000000000";
      when "010001100001011" => color_data <= "000000000000";
      when "010001100001100" => color_data <= "000000000000";
      when "010001100001101" => color_data <= "000000000000";
      when "010001100001110" => color_data <= "000000000000";
      when "010001100001111" => color_data <= "000000000000";
      when "010001100010000" => color_data <= "000000000000";
      when "010001100010001" => color_data <= "000000000000";
      when "010001100010010" => color_data <= "000000000000";
      when "010001100010011" => color_data <= "000000000000";
      when "010001100010100" => color_data <= "000000000000";
      when "010001100010101" => color_data <= "000000000000";
      when "010001100010110" => color_data <= "000000000000";
      when "010001100010111" => color_data <= "000000000000";
      when "010001100011000" => color_data <= "100001110010";
      when "010001100011001" => color_data <= "110110100000";
      when "010001100011010" => color_data <= "111111000001";
      when "010001100011011" => color_data <= "110110100000";
      when "010001100011100" => color_data <= "010101010011";
      when "010001100011101" => color_data <= "000000000000";
      when "010001100011110" => color_data <= "000000000000";
      when "010001100011111" => color_data <= "000000000000";
      when "010001100100000" => color_data <= "000000000000";
      when "010001100100001" => color_data <= "000000000000";
      when "010001100100010" => color_data <= "000000000000";
      when "010001100100011" => color_data <= "000000000000";
      when "010001100100100" => color_data <= "000000000000";
      when "010001100100101" => color_data <= "000000000000";
      when "010001100100110" => color_data <= "000000000000";
      when "010001100100111" => color_data <= "000000000000";
      when "010001100101000" => color_data <= "000000000000";
      when "010001100101001" => color_data <= "000000000000";
      when "010001100101010" => color_data <= "000000000000";
      when "010001100101011" => color_data <= "000000000000";
      when "010001100101100" => color_data <= "000000000000";
      when "010001100101101" => color_data <= "000000000000";
      when "010001100101110" => color_data <= "000000000000";
      when "010001100101111" => color_data <= "000000000000";
      when "010001100110000" => color_data <= "000000000000";
      when "010001100110001" => color_data <= "000000000000";
      when "010001100110010" => color_data <= "000000000000";
      when "010001100110011" => color_data <= "000000000000";
      when "010001100110100" => color_data <= "000000000000";
      when "010001100110101" => color_data <= "000000000000";
      when "010001100110110" => color_data <= "000000000000";
      when "010001100110111" => color_data <= "000000000000";
      when "010001100111000" => color_data <= "000000000000";
      when "010001100111001" => color_data <= "000000000000";
      when "010001100111010" => color_data <= "000000000000";
      when "010001100111011" => color_data <= "000000000000";
      when "010001100111100" => color_data <= "000000000000";
      when "010001100111101" => color_data <= "000000000000";
      when "010001100111110" => color_data <= "000000000000";
      when "010001100111111" => color_data <= "000000000000";
      when "010001101000000" => color_data <= "000000000000";
      when "010001101000001" => color_data <= "000000000000";
      when "010001101000010" => color_data <= "000000000000";
      when "010001101000011" => color_data <= "000000000000";
      when "010001101000100" => color_data <= "000000000000";
      when "010001101000101" => color_data <= "000000000000";
      when "010001101000110" => color_data <= "000000000000";
      when "010001101000111" => color_data <= "000000000000";
      when "010001101001000" => color_data <= "000000000000";
      when "010001101001001" => color_data <= "000000000000";
      when "010001101001010" => color_data <= "000000000000";
      when "010001101001011" => color_data <= "110010010001";
      when "010001101001100" => color_data <= "111110110000";
      when "010001101001101" => color_data <= "111111000000";
      when "010001101001110" => color_data <= "110110100000";
      when "010001101001111" => color_data <= "000100010001";
      when "010001101010000" => color_data <= "000000000000";
      when "010001101010001" => color_data <= "000000000000";
      when "010001101010010" => color_data <= "000000000000";
      when "010001101010011" => color_data <= "000000000000";
      when "010001101010100" => color_data <= "000000000000";
      when "010001101010101" => color_data <= "000000000000";
      when "010001101010110" => color_data <= "000000000000";
      when "010001101010111" => color_data <= "000000000000";
      when "010001101011000" => color_data <= "000000000000";
      when "010001101011001" => color_data <= "000000000000";
      when "010001101011010" => color_data <= "000000000000";
      when "010001101011011" => color_data <= "000000000000";
      when "010001101011100" => color_data <= "000000000000";
      when "010001101011101" => color_data <= "000000000000";
      when "010001101011110" => color_data <= "000000000000";
      when "010001101011111" => color_data <= "000000000000";
      when "010001101100000" => color_data <= "000000000000";
      when "010001101100001" => color_data <= "000000000000";
      when "010001101100010" => color_data <= "000000000000";
      when "010001101100011" => color_data <= "000000000000";
      when "010001110000000" => color_data <= "000000000000";
      when "010001110000001" => color_data <= "000000000000";
      when "010001110000010" => color_data <= "000000000000";
      when "010001110000011" => color_data <= "000000000000";
      when "010001110000100" => color_data <= "000000000000";
      when "010001110000101" => color_data <= "000000000000";
      when "010001110000110" => color_data <= "000000000000";
      when "010001110000111" => color_data <= "000000000000";
      when "010001110001000" => color_data <= "000000000000";
      when "010001110001001" => color_data <= "000000000000";
      when "010001110001010" => color_data <= "000000000000";
      when "010001110001011" => color_data <= "000000000000";
      when "010001110001100" => color_data <= "000000000000";
      when "010001110001101" => color_data <= "000000000000";
      when "010001110001110" => color_data <= "000000000000";
      when "010001110001111" => color_data <= "000000000000";
      when "010001110010000" => color_data <= "000000000000";
      when "010001110010001" => color_data <= "000000000000";
      when "010001110010010" => color_data <= "000000000000";
      when "010001110010011" => color_data <= "000000000000";
      when "010001110010100" => color_data <= "000000000000";
      when "010001110010101" => color_data <= "000000000000";
      when "010001110010110" => color_data <= "000000000000";
      when "010001110010111" => color_data <= "000000000000";
      when "010001110011000" => color_data <= "000000000000";
      when "010001110011001" => color_data <= "101010000010";
      when "010001110011010" => color_data <= "110110100000";
      when "010001110011011" => color_data <= "111111000000";
      when "010001110011100" => color_data <= "110110100000";
      when "010001110011101" => color_data <= "001100110010";
      when "010001110011110" => color_data <= "000000000000";
      when "010001110011111" => color_data <= "000000000000";
      when "010001110100000" => color_data <= "000000000000";
      when "010001110100001" => color_data <= "000000000000";
      when "010001110100010" => color_data <= "000000000000";
      when "010001110100011" => color_data <= "000000000000";
      when "010001110100100" => color_data <= "000000000000";
      when "010001110100101" => color_data <= "000000000000";
      when "010001110100110" => color_data <= "000000000000";
      when "010001110100111" => color_data <= "000000000000";
      when "010001110101000" => color_data <= "000000000000";
      when "010001110101001" => color_data <= "000000000000";
      when "010001110101010" => color_data <= "000000000000";
      when "010001110101011" => color_data <= "000000000000";
      when "010001110101100" => color_data <= "000000000000";
      when "010001110101101" => color_data <= "000000000000";
      when "010001110101110" => color_data <= "000000000000";
      when "010001110101111" => color_data <= "000000000000";
      when "010001110110000" => color_data <= "000000000000";
      when "010001110110001" => color_data <= "000000000000";
      when "010001110110010" => color_data <= "000000000000";
      when "010001110110011" => color_data <= "000000000000";
      when "010001110110100" => color_data <= "000000000000";
      when "010001110110101" => color_data <= "000000000000";
      when "010001110110110" => color_data <= "000000000000";
      when "010001110110111" => color_data <= "000000000000";
      when "010001110111000" => color_data <= "000000000000";
      when "010001110111001" => color_data <= "000000000000";
      when "010001110111010" => color_data <= "000000000000";
      when "010001110111011" => color_data <= "000000000000";
      when "010001110111100" => color_data <= "000000000000";
      when "010001110111101" => color_data <= "000000000000";
      when "010001110111110" => color_data <= "000000000000";
      when "010001110111111" => color_data <= "000000000000";
      when "010001111000000" => color_data <= "000000000000";
      when "010001111000001" => color_data <= "000000000000";
      when "010001111000010" => color_data <= "000000000000";
      when "010001111000011" => color_data <= "000000000000";
      when "010001111000100" => color_data <= "000000000000";
      when "010001111000101" => color_data <= "000000000000";
      when "010001111000110" => color_data <= "000000000000";
      when "010001111000111" => color_data <= "000000000000";
      when "010001111001000" => color_data <= "000000000000";
      when "010001111001001" => color_data <= "000000000000";
      when "010001111001010" => color_data <= "101110010001";
      when "010001111001011" => color_data <= "110110100000";
      when "010001111001100" => color_data <= "111111000000";
      when "010001111001101" => color_data <= "110110100000";
      when "010001111001110" => color_data <= "001100110010";
      when "010001111001111" => color_data <= "000000000000";
      when "010001111010000" => color_data <= "000000000000";
      when "010001111010001" => color_data <= "000000000000";
      when "010001111010010" => color_data <= "000000000000";
      when "010001111010011" => color_data <= "000000000000";
      when "010001111010100" => color_data <= "000000000000";
      when "010001111010101" => color_data <= "000000000000";
      when "010001111010110" => color_data <= "000000000000";
      when "010001111010111" => color_data <= "000000000000";
      when "010001111011000" => color_data <= "000000000000";
      when "010001111011001" => color_data <= "000000000000";
      when "010001111011010" => color_data <= "000000000000";
      when "010001111011011" => color_data <= "000000000000";
      when "010001111011100" => color_data <= "000000000000";
      when "010001111011101" => color_data <= "000000000000";
      when "010001111011110" => color_data <= "000000000000";
      when "010001111011111" => color_data <= "000000000000";
      when "010001111100000" => color_data <= "000000000000";
      when "010001111100001" => color_data <= "000000000000";
      when "010001111100010" => color_data <= "000000000000";
      when "010001111100011" => color_data <= "000000000000";
      when "010010000000000" => color_data <= "000000000000";
      when "010010000000001" => color_data <= "000000000000";
      when "010010000000010" => color_data <= "000000000000";
      when "010010000000011" => color_data <= "000000000000";
      when "010010000000100" => color_data <= "000000000000";
      when "010010000000101" => color_data <= "000000000000";
      when "010010000000110" => color_data <= "000000000000";
      when "010010000000111" => color_data <= "000000000000";
      when "010010000001000" => color_data <= "000000000000";
      when "010010000001001" => color_data <= "000000000000";
      when "010010000001010" => color_data <= "000000000000";
      when "010010000001011" => color_data <= "000000000000";
      when "010010000001100" => color_data <= "000000000000";
      when "010010000001101" => color_data <= "000000000000";
      when "010010000001110" => color_data <= "000000000000";
      when "010010000001111" => color_data <= "000000000000";
      when "010010000010000" => color_data <= "000000000000";
      when "010010000010001" => color_data <= "000000000000";
      when "010010000010010" => color_data <= "000000000000";
      when "010010000010011" => color_data <= "000000000000";
      when "010010000010100" => color_data <= "000000000000";
      when "010010000010101" => color_data <= "000000000000";
      when "010010000010110" => color_data <= "000000000000";
      when "010010000010111" => color_data <= "000000000000";
      when "010010000011000" => color_data <= "000000000000";
      when "010010000011001" => color_data <= "000000000000";
      when "010010000011010" => color_data <= "110010010001";
      when "010010000011011" => color_data <= "111110110000";
      when "010010000011100" => color_data <= "111111000000";
      when "010010000011101" => color_data <= "110110100000";
      when "010010000011110" => color_data <= "001000100001";
      when "010010000011111" => color_data <= "000000000000";
      when "010010000100000" => color_data <= "000000000000";
      when "010010000100001" => color_data <= "000000000000";
      when "010010000100010" => color_data <= "000000000000";
      when "010010000100011" => color_data <= "000000000000";
      when "010010000100100" => color_data <= "000000000000";
      when "010010000100101" => color_data <= "000000000000";
      when "010010000100110" => color_data <= "000000000000";
      when "010010000100111" => color_data <= "000000000000";
      when "010010000101000" => color_data <= "000000000000";
      when "010010000101001" => color_data <= "000000000000";
      when "010010000101010" => color_data <= "000000000000";
      when "010010000101011" => color_data <= "000000000000";
      when "010010000101100" => color_data <= "000000000000";
      when "010010000101101" => color_data <= "000000000000";
      when "010010000101110" => color_data <= "000000000000";
      when "010010000101111" => color_data <= "000000000000";
      when "010010000110000" => color_data <= "000000000000";
      when "010010000110001" => color_data <= "000000000000";
      when "010010000110010" => color_data <= "000000000000";
      when "010010000110011" => color_data <= "000000000000";
      when "010010000110100" => color_data <= "000000000000";
      when "010010000110101" => color_data <= "000000000000";
      when "010010000110110" => color_data <= "000000000000";
      when "010010000110111" => color_data <= "000000000000";
      when "010010000111000" => color_data <= "000000000000";
      when "010010000111001" => color_data <= "000000000000";
      when "010010000111010" => color_data <= "000000000000";
      when "010010000111011" => color_data <= "000000000000";
      when "010010000111100" => color_data <= "000000000000";
      when "010010000111101" => color_data <= "000000000000";
      when "010010000111110" => color_data <= "000000000000";
      when "010010000111111" => color_data <= "000000000000";
      when "010010001000000" => color_data <= "000000000000";
      when "010010001000001" => color_data <= "000000000000";
      when "010010001000010" => color_data <= "000000000000";
      when "010010001000011" => color_data <= "000000000000";
      when "010010001000100" => color_data <= "000000000000";
      when "010010001000101" => color_data <= "000000000000";
      when "010010001000110" => color_data <= "000000000000";
      when "010010001000111" => color_data <= "000000000000";
      when "010010001001000" => color_data <= "000000000000";
      when "010010001001001" => color_data <= "101010000010";
      when "010010001001010" => color_data <= "110110100000";
      when "010010001001011" => color_data <= "111111000000";
      when "010010001001100" => color_data <= "110110100000";
      when "010010001001101" => color_data <= "010001000010";
      when "010010001001110" => color_data <= "000000000000";
      when "010010001001111" => color_data <= "000000000000";
      when "010010001010000" => color_data <= "000000000000";
      when "010010001010001" => color_data <= "000000000000";
      when "010010001010010" => color_data <= "000000000000";
      when "010010001010011" => color_data <= "000000000000";
      when "010010001010100" => color_data <= "000000000000";
      when "010010001010101" => color_data <= "000000000000";
      when "010010001010110" => color_data <= "000000000000";
      when "010010001010111" => color_data <= "000000000000";
      when "010010001011000" => color_data <= "000000000000";
      when "010010001011001" => color_data <= "000000000000";
      when "010010001011010" => color_data <= "000000000000";
      when "010010001011011" => color_data <= "000000000000";
      when "010010001011100" => color_data <= "000000000000";
      when "010010001011101" => color_data <= "000000000000";
      when "010010001011110" => color_data <= "000000000000";
      when "010010001011111" => color_data <= "000000000000";
      when "010010001100000" => color_data <= "000000000000";
      when "010010001100001" => color_data <= "000000000000";
      when "010010001100010" => color_data <= "000000000000";
      when "010010001100011" => color_data <= "000000000000";
      when "010010010000000" => color_data <= "000000000000";
      when "010010010000001" => color_data <= "000000000000";
      when "010010010000010" => color_data <= "000000000000";
      when "010010010000011" => color_data <= "000000000000";
      when "010010010000100" => color_data <= "000000000000";
      when "010010010000101" => color_data <= "000000000000";
      when "010010010000110" => color_data <= "000000000000";
      when "010010010000111" => color_data <= "000000000000";
      when "010010010001000" => color_data <= "000000000000";
      when "010010010001001" => color_data <= "000000000000";
      when "010010010001010" => color_data <= "000000000000";
      when "010010010001011" => color_data <= "000000000000";
      when "010010010001100" => color_data <= "000000000000";
      when "010010010001101" => color_data <= "000000000000";
      when "010010010001110" => color_data <= "000000000000";
      when "010010010001111" => color_data <= "000000000000";
      when "010010010010000" => color_data <= "000000000000";
      when "010010010010001" => color_data <= "000000000000";
      when "010010010010010" => color_data <= "000000000000";
      when "010010010010011" => color_data <= "000000000000";
      when "010010010010100" => color_data <= "000000000000";
      when "010010010010101" => color_data <= "000000000000";
      when "010010010010110" => color_data <= "000000000000";
      when "010010010010111" => color_data <= "000000000000";
      when "010010010011000" => color_data <= "000000000000";
      when "010010010011001" => color_data <= "000000000000";
      when "010010010011010" => color_data <= "000000000000";
      when "010010010011011" => color_data <= "110010010000";
      when "010010010011100" => color_data <= "111110110000";
      when "010010010011101" => color_data <= "111110110000";
      when "010010010011110" => color_data <= "110110100000";
      when "010010010011111" => color_data <= "000100010001";
      when "010010010100000" => color_data <= "000000000000";
      when "010010010100001" => color_data <= "000000000000";
      when "010010010100010" => color_data <= "000000000000";
      when "010010010100011" => color_data <= "000000000000";
      when "010010010100100" => color_data <= "000000000000";
      when "010010010100101" => color_data <= "000000000000";
      when "010010010100110" => color_data <= "000000000000";
      when "010010010100111" => color_data <= "000000000000";
      when "010010010101000" => color_data <= "000000000000";
      when "010010010101001" => color_data <= "000000000000";
      when "010010010101010" => color_data <= "000000000000";
      when "010010010101011" => color_data <= "000000000000";
      when "010010010101100" => color_data <= "000000000000";
      when "010010010101101" => color_data <= "000000000000";
      when "010010010101110" => color_data <= "000000000000";
      when "010010010101111" => color_data <= "000000000000";
      when "010010010110000" => color_data <= "000000000000";
      when "010010010110001" => color_data <= "000000000000";
      when "010010010110010" => color_data <= "000000000000";
      when "010010010110011" => color_data <= "000000000000";
      when "010010010110100" => color_data <= "000000000000";
      when "010010010110101" => color_data <= "000000000000";
      when "010010010110110" => color_data <= "000000000000";
      when "010010010110111" => color_data <= "000000000000";
      when "010010010111000" => color_data <= "000000000000";
      when "010010010111001" => color_data <= "000000000000";
      when "010010010111010" => color_data <= "000000000000";
      when "010010010111011" => color_data <= "000000000000";
      when "010010010111100" => color_data <= "000000000000";
      when "010010010111101" => color_data <= "000000000000";
      when "010010010111110" => color_data <= "000000000000";
      when "010010010111111" => color_data <= "000000000000";
      when "010010011000000" => color_data <= "000000000000";
      when "010010011000001" => color_data <= "000000000000";
      when "010010011000010" => color_data <= "000000000000";
      when "010010011000011" => color_data <= "000000000000";
      when "010010011000100" => color_data <= "000000000000";
      when "010010011000101" => color_data <= "000000000000";
      when "010010011000110" => color_data <= "000000000000";
      when "010010011000111" => color_data <= "000000000000";
      when "010010011001000" => color_data <= "101010000010";
      when "010010011001001" => color_data <= "110110100000";
      when "010010011001010" => color_data <= "111111000000";
      when "010010011001011" => color_data <= "110110100000";
      when "010010011001100" => color_data <= "010101010010";
      when "010010011001101" => color_data <= "000000000000";
      when "010010011001110" => color_data <= "000000000000";
      when "010010011001111" => color_data <= "000000000000";
      when "010010011010000" => color_data <= "000000000000";
      when "010010011010001" => color_data <= "000000000000";
      when "010010011010010" => color_data <= "000000000000";
      when "010010011010011" => color_data <= "000000000000";
      when "010010011010100" => color_data <= "000000000000";
      when "010010011010101" => color_data <= "000000000000";
      when "010010011010110" => color_data <= "000000000000";
      when "010010011010111" => color_data <= "000000000000";
      when "010010011011000" => color_data <= "000000000000";
      when "010010011011001" => color_data <= "000000000000";
      when "010010011011010" => color_data <= "000000000000";
      when "010010011011011" => color_data <= "000000000000";
      when "010010011011100" => color_data <= "000000000000";
      when "010010011011101" => color_data <= "000000000000";
      when "010010011011110" => color_data <= "000000000000";
      when "010010011011111" => color_data <= "000000000000";
      when "010010011100000" => color_data <= "000000000000";
      when "010010011100001" => color_data <= "000000000000";
      when "010010011100010" => color_data <= "000000000000";
      when "010010011100011" => color_data <= "000000000000";
      when "010010100000000" => color_data <= "000000000000";
      when "010010100000001" => color_data <= "000000000000";
      when "010010100000010" => color_data <= "000000000000";
      when "010010100000011" => color_data <= "000000000000";
      when "010010100000100" => color_data <= "000000000000";
      when "010010100000101" => color_data <= "000000000000";
      when "010010100000110" => color_data <= "000000000000";
      when "010010100000111" => color_data <= "000000000000";
      when "010010100001000" => color_data <= "000000000000";
      when "010010100001001" => color_data <= "000000000000";
      when "010010100001010" => color_data <= "000000000000";
      when "010010100001011" => color_data <= "000000000000";
      when "010010100001100" => color_data <= "000000000000";
      when "010010100001101" => color_data <= "000000000000";
      when "010010100001110" => color_data <= "000000000000";
      when "010010100001111" => color_data <= "000000000000";
      when "010010100010000" => color_data <= "000000000000";
      when "010010100010001" => color_data <= "000000000000";
      when "010010100010010" => color_data <= "000000000000";
      when "010010100010011" => color_data <= "000000000000";
      when "010010100010100" => color_data <= "000000000000";
      when "010010100010101" => color_data <= "000000000000";
      when "010010100010110" => color_data <= "000000000000";
      when "010010100010111" => color_data <= "000000000000";
      when "010010100011000" => color_data <= "000000000000";
      when "010010100011001" => color_data <= "000000000000";
      when "010010100011010" => color_data <= "000000000000";
      when "010010100011011" => color_data <= "000000000000";
      when "010010100011100" => color_data <= "110110100000";
      when "010010100011101" => color_data <= "111111000000";
      when "010010100011110" => color_data <= "111110110000";
      when "010010100011111" => color_data <= "110110010000";
      when "010010100100000" => color_data <= "000100010001";
      when "010010100100001" => color_data <= "000000000000";
      when "010010100100010" => color_data <= "000000000000";
      when "010010100100011" => color_data <= "000000000000";
      when "010010100100100" => color_data <= "000000000000";
      when "010010100100101" => color_data <= "000000000000";
      when "010010100100110" => color_data <= "000000000000";
      when "010010100100111" => color_data <= "000000000000";
      when "010010100101000" => color_data <= "000000000000";
      when "010010100101001" => color_data <= "000000000000";
      when "010010100101010" => color_data <= "000000000000";
      when "010010100101011" => color_data <= "000000000000";
      when "010010100101100" => color_data <= "000000000000";
      when "010010100101101" => color_data <= "000000000000";
      when "010010100101110" => color_data <= "000000000000";
      when "010010100101111" => color_data <= "000000000000";
      when "010010100110000" => color_data <= "000000000000";
      when "010010100110001" => color_data <= "000000000000";
      when "010010100110010" => color_data <= "000000000000";
      when "010010100110011" => color_data <= "000000000000";
      when "010010100110100" => color_data <= "000000000000";
      when "010010100110101" => color_data <= "000000000000";
      when "010010100110110" => color_data <= "000000000000";
      when "010010100110111" => color_data <= "000000000000";
      when "010010100111000" => color_data <= "000000000000";
      when "010010100111001" => color_data <= "000000000000";
      when "010010100111010" => color_data <= "000000000000";
      when "010010100111011" => color_data <= "000000000000";
      when "010010100111100" => color_data <= "000000000000";
      when "010010100111101" => color_data <= "000000000000";
      when "010010100111110" => color_data <= "000000000000";
      when "010010100111111" => color_data <= "000000000000";
      when "010010101000000" => color_data <= "000000000000";
      when "010010101000001" => color_data <= "000000000000";
      when "010010101000010" => color_data <= "000000000000";
      when "010010101000011" => color_data <= "000000000000";
      when "010010101000100" => color_data <= "000000000000";
      when "010010101000101" => color_data <= "000000000000";
      when "010010101000110" => color_data <= "000000000000";
      when "010010101000111" => color_data <= "101010000010";
      when "010010101001000" => color_data <= "110110100000";
      when "010010101001001" => color_data <= "111111000000";
      when "010010101001010" => color_data <= "110110100000";
      when "010010101001011" => color_data <= "010101010011";
      when "010010101001100" => color_data <= "000000000000";
      when "010010101001101" => color_data <= "000000000000";
      when "010010101001110" => color_data <= "000000000000";
      when "010010101001111" => color_data <= "000000000000";
      when "010010101010000" => color_data <= "000000000000";
      when "010010101010001" => color_data <= "000000000000";
      when "010010101010010" => color_data <= "000000000000";
      when "010010101010011" => color_data <= "000000000000";
      when "010010101010100" => color_data <= "000000000000";
      when "010010101010101" => color_data <= "000000000000";
      when "010010101010110" => color_data <= "000000000000";
      when "010010101010111" => color_data <= "000000000000";
      when "010010101011000" => color_data <= "000000000000";
      when "010010101011001" => color_data <= "000000000000";
      when "010010101011010" => color_data <= "000000000000";
      when "010010101011011" => color_data <= "000000000000";
      when "010010101011100" => color_data <= "000000000000";
      when "010010101011101" => color_data <= "000000000000";
      when "010010101011110" => color_data <= "000000000000";
      when "010010101011111" => color_data <= "000000000000";
      when "010010101100000" => color_data <= "000000000000";
      when "010010101100001" => color_data <= "000000000000";
      when "010010101100010" => color_data <= "000000000000";
      when "010010101100011" => color_data <= "000000000000";
      when "010010110000000" => color_data <= "000000000000";
      when "010010110000001" => color_data <= "000000000000";
      when "010010110000010" => color_data <= "000000000000";
      when "010010110000011" => color_data <= "000000000000";
      when "010010110000100" => color_data <= "000000000000";
      when "010010110000101" => color_data <= "000000000000";
      when "010010110000110" => color_data <= "000000000000";
      when "010010110000111" => color_data <= "000000000000";
      when "010010110001000" => color_data <= "000000000000";
      when "010010110001001" => color_data <= "000000000000";
      when "010010110001010" => color_data <= "000000000000";
      when "010010110001011" => color_data <= "000000000000";
      when "010010110001100" => color_data <= "000000000000";
      when "010010110001101" => color_data <= "000000000000";
      when "010010110001110" => color_data <= "000000000000";
      when "010010110001111" => color_data <= "000000000000";
      when "010010110010000" => color_data <= "000000000000";
      when "010010110010001" => color_data <= "000000000000";
      when "010010110010010" => color_data <= "000000000000";
      when "010010110010011" => color_data <= "000000000000";
      when "010010110010100" => color_data <= "000000000000";
      when "010010110010101" => color_data <= "000000000000";
      when "010010110010110" => color_data <= "000000000000";
      when "010010110010111" => color_data <= "000000000000";
      when "010010110011000" => color_data <= "000000000000";
      when "010010110011001" => color_data <= "000000000000";
      when "010010110011010" => color_data <= "000000000000";
      when "010010110011011" => color_data <= "000000000000";
      when "010010110011100" => color_data <= "000000000000";
      when "010010110011101" => color_data <= "110010010000";
      when "010010110011110" => color_data <= "111110110000";
      when "010010110011111" => color_data <= "111110110000";
      when "010010110100000" => color_data <= "110110100000";
      when "010010110100001" => color_data <= "000100010001";
      when "010010110100010" => color_data <= "000000000000";
      when "010010110100011" => color_data <= "000000000000";
      when "010010110100100" => color_data <= "000000000000";
      when "010010110100101" => color_data <= "000000000000";
      when "010010110100110" => color_data <= "000000000000";
      when "010010110100111" => color_data <= "000000000000";
      when "010010110101000" => color_data <= "000000000000";
      when "010010110101001" => color_data <= "000000000000";
      when "010010110101010" => color_data <= "000000000000";
      when "010010110101011" => color_data <= "000000000000";
      when "010010110101100" => color_data <= "000000000000";
      when "010010110101101" => color_data <= "000000000000";
      when "010010110101110" => color_data <= "000000000000";
      when "010010110101111" => color_data <= "000000000000";
      when "010010110110000" => color_data <= "000000000000";
      when "010010110110001" => color_data <= "000000000000";
      when "010010110110010" => color_data <= "000000000000";
      when "010010110110011" => color_data <= "000000000000";
      when "010010110110100" => color_data <= "000000000000";
      when "010010110110101" => color_data <= "000000000000";
      when "010010110110110" => color_data <= "000000000000";
      when "010010110110111" => color_data <= "000000000000";
      when "010010110111000" => color_data <= "000000000000";
      when "010010110111001" => color_data <= "000000000000";
      when "010010110111010" => color_data <= "000000000000";
      when "010010110111011" => color_data <= "000000000000";
      when "010010110111100" => color_data <= "000000000000";
      when "010010110111101" => color_data <= "000000000000";
      when "010010110111110" => color_data <= "000000000000";
      when "010010110111111" => color_data <= "000000000000";
      when "010010111000000" => color_data <= "000000000000";
      when "010010111000001" => color_data <= "000000000000";
      when "010010111000010" => color_data <= "000000000000";
      when "010010111000011" => color_data <= "000000000000";
      when "010010111000100" => color_data <= "000000000000";
      when "010010111000101" => color_data <= "000000000000";
      when "010010111000110" => color_data <= "101010000010";
      when "010010111000111" => color_data <= "110110100000";
      when "010010111001000" => color_data <= "111111000000";
      when "010010111001001" => color_data <= "110110100000";
      when "010010111001010" => color_data <= "010101000010";
      when "010010111001011" => color_data <= "000000000000";
      when "010010111001100" => color_data <= "000000000000";
      when "010010111001101" => color_data <= "000000000000";
      when "010010111001110" => color_data <= "000000000000";
      when "010010111001111" => color_data <= "000000000000";
      when "010010111010000" => color_data <= "000000000000";
      when "010010111010001" => color_data <= "000000000000";
      when "010010111010010" => color_data <= "000000000000";
      when "010010111010011" => color_data <= "000000000000";
      when "010010111010100" => color_data <= "000000000000";
      when "010010111010101" => color_data <= "000000000000";
      when "010010111010110" => color_data <= "000000000000";
      when "010010111010111" => color_data <= "000000000000";
      when "010010111011000" => color_data <= "000000000000";
      when "010010111011001" => color_data <= "000000000000";
      when "010010111011010" => color_data <= "000000000000";
      when "010010111011011" => color_data <= "000000000000";
      when "010010111011100" => color_data <= "000000000000";
      when "010010111011101" => color_data <= "000000000000";
      when "010010111011110" => color_data <= "000000000000";
      when "010010111011111" => color_data <= "000000000000";
      when "010010111100000" => color_data <= "000000000000";
      when "010010111100001" => color_data <= "000000000000";
      when "010010111100010" => color_data <= "000000000000";
      when "010010111100011" => color_data <= "000000000000";
      when "010011000000000" => color_data <= "000000000000";
      when "010011000000001" => color_data <= "000000000000";
      when "010011000000010" => color_data <= "000000000000";
      when "010011000000011" => color_data <= "000000000000";
      when "010011000000100" => color_data <= "000000000000";
      when "010011000000101" => color_data <= "000000000000";
      when "010011000000110" => color_data <= "000000000000";
      when "010011000000111" => color_data <= "000000000000";
      when "010011000001000" => color_data <= "000000000000";
      when "010011000001001" => color_data <= "000000000000";
      when "010011000001010" => color_data <= "000000000000";
      when "010011000001011" => color_data <= "000000000000";
      when "010011000001100" => color_data <= "000000000000";
      when "010011000001101" => color_data <= "000000000000";
      when "010011000001110" => color_data <= "000000000000";
      when "010011000001111" => color_data <= "000000000000";
      when "010011000010000" => color_data <= "000000000000";
      when "010011000010001" => color_data <= "000000000000";
      when "010011000010010" => color_data <= "000000000000";
      when "010011000010011" => color_data <= "000000000000";
      when "010011000010100" => color_data <= "000000000000";
      when "010011000010101" => color_data <= "000000000000";
      when "010011000010110" => color_data <= "000000000000";
      when "010011000010111" => color_data <= "000000000000";
      when "010011000011000" => color_data <= "000000000000";
      when "010011000011001" => color_data <= "000000000000";
      when "010011000011010" => color_data <= "000000000000";
      when "010011000011011" => color_data <= "000000000000";
      when "010011000011100" => color_data <= "000000000000";
      when "010011000011101" => color_data <= "000000000000";
      when "010011000011110" => color_data <= "110010010000";
      when "010011000011111" => color_data <= "110110100000";
      when "010011000100000" => color_data <= "111110110000";
      when "010011000100001" => color_data <= "110010010001";
      when "010011000100010" => color_data <= "000100010001";
      when "010011000100011" => color_data <= "000000000000";
      when "010011000100100" => color_data <= "000000000000";
      when "010011000100101" => color_data <= "000000000000";
      when "010011000100110" => color_data <= "000000000000";
      when "010011000100111" => color_data <= "000000000000";
      when "010011000101000" => color_data <= "000000000000";
      when "010011000101001" => color_data <= "000000000000";
      when "010011000101010" => color_data <= "000000000000";
      when "010011000101011" => color_data <= "000000000000";
      when "010011000101100" => color_data <= "000000000000";
      when "010011000101101" => color_data <= "000000000000";
      when "010011000101110" => color_data <= "000000000000";
      when "010011000101111" => color_data <= "000000000000";
      when "010011000110000" => color_data <= "000000000000";
      when "010011000110001" => color_data <= "000000000000";
      when "010011000110010" => color_data <= "000000000000";
      when "010011000110011" => color_data <= "000000000000";
      when "010011000110100" => color_data <= "000000000000";
      when "010011000110101" => color_data <= "000000000000";
      when "010011000110110" => color_data <= "000000000000";
      when "010011000110111" => color_data <= "000000000000";
      when "010011000111000" => color_data <= "000000000000";
      when "010011000111001" => color_data <= "000000000000";
      when "010011000111010" => color_data <= "000000000000";
      when "010011000111011" => color_data <= "000000000000";
      when "010011000111100" => color_data <= "000000000000";
      when "010011000111101" => color_data <= "000000000000";
      when "010011000111110" => color_data <= "000000000000";
      when "010011000111111" => color_data <= "000000000000";
      when "010011001000000" => color_data <= "000000000000";
      when "010011001000001" => color_data <= "000000000000";
      when "010011001000010" => color_data <= "000000000000";
      when "010011001000011" => color_data <= "000000000000";
      when "010011001000100" => color_data <= "000000000000";
      when "010011001000101" => color_data <= "101010000001";
      when "010011001000110" => color_data <= "110110100000";
      when "010011001000111" => color_data <= "111111000000";
      when "010011001001000" => color_data <= "110110100000";
      when "010011001001001" => color_data <= "010001000010";
      when "010011001001010" => color_data <= "000000000000";
      when "010011001001011" => color_data <= "000000000000";
      when "010011001001100" => color_data <= "000000000000";
      when "010011001001101" => color_data <= "000000000000";
      when "010011001001110" => color_data <= "000000000000";
      when "010011001001111" => color_data <= "000000000000";
      when "010011001010000" => color_data <= "000000000000";
      when "010011001010001" => color_data <= "000000000000";
      when "010011001010010" => color_data <= "000000000000";
      when "010011001010011" => color_data <= "000000000000";
      when "010011001010100" => color_data <= "000000000000";
      when "010011001010101" => color_data <= "000000000000";
      when "010011001010110" => color_data <= "000000000000";
      when "010011001010111" => color_data <= "000000000000";
      when "010011001011000" => color_data <= "000000000000";
      when "010011001011001" => color_data <= "000000000000";
      when "010011001011010" => color_data <= "000000000000";
      when "010011001011011" => color_data <= "000000000000";
      when "010011001011100" => color_data <= "000000000000";
      when "010011001011101" => color_data <= "000000000000";
      when "010011001011110" => color_data <= "000000000000";
      when "010011001011111" => color_data <= "000000000000";
      when "010011001100000" => color_data <= "000000000000";
      when "010011001100001" => color_data <= "000000000000";
      when "010011001100010" => color_data <= "000000000000";
      when "010011001100011" => color_data <= "000000000000";
      when "010011010000000" => color_data <= "000000000000";
      when "010011010000001" => color_data <= "000000000000";
      when "010011010000010" => color_data <= "000000000000";
      when "010011010000011" => color_data <= "000000000000";
      when "010011010000100" => color_data <= "000000000000";
      when "010011010000101" => color_data <= "000000000000";
      when "010011010000110" => color_data <= "000000000000";
      when "010011010000111" => color_data <= "000000000000";
      when "010011010001000" => color_data <= "000000000000";
      when "010011010001001" => color_data <= "000000000000";
      when "010011010001010" => color_data <= "000000000000";
      when "010011010001011" => color_data <= "000000000000";
      when "010011010001100" => color_data <= "000000000000";
      when "010011010001101" => color_data <= "000000000000";
      when "010011010001110" => color_data <= "000000000000";
      when "010011010001111" => color_data <= "000000000000";
      when "010011010010000" => color_data <= "000000000000";
      when "010011010010001" => color_data <= "000000000000";
      when "010011010010010" => color_data <= "000000000000";
      when "010011010010011" => color_data <= "000000000000";
      when "010011010010100" => color_data <= "000000000000";
      when "010011010010101" => color_data <= "000000000000";
      when "010011010010110" => color_data <= "000000000000";
      when "010011010010111" => color_data <= "000000000000";
      when "010011010011000" => color_data <= "000000000000";
      when "010011010011001" => color_data <= "000000000000";
      when "010011010011010" => color_data <= "000000000000";
      when "010011010011011" => color_data <= "000000000000";
      when "010011010011100" => color_data <= "000000000000";
      when "010011010011101" => color_data <= "000000000000";
      when "010011010011110" => color_data <= "000000000000";
      when "010011010011111" => color_data <= "101010000001";
      when "010011010100000" => color_data <= "110110100000";
      when "010011010100001" => color_data <= "111110110000";
      when "010011010100010" => color_data <= "110110100000";
      when "010011010100011" => color_data <= "001100110010";
      when "010011010100100" => color_data <= "000000000000";
      when "010011010100101" => color_data <= "000000000000";
      when "010011010100110" => color_data <= "000000000000";
      when "010011010100111" => color_data <= "000000000000";
      when "010011010101000" => color_data <= "000000000000";
      when "010011010101001" => color_data <= "000000000000";
      when "010011010101010" => color_data <= "000000000000";
      when "010011010101011" => color_data <= "000000000000";
      when "010011010101100" => color_data <= "000000000000";
      when "010011010101101" => color_data <= "000000000000";
      when "010011010101110" => color_data <= "000000000000";
      when "010011010101111" => color_data <= "000000000000";
      when "010011010110000" => color_data <= "000000000000";
      when "010011010110001" => color_data <= "000000000000";
      when "010011010110010" => color_data <= "000000000000";
      when "010011010110011" => color_data <= "000000000000";
      when "010011010110100" => color_data <= "000000000000";
      when "010011010110101" => color_data <= "000000000000";
      when "010011010110110" => color_data <= "000000000000";
      when "010011010110111" => color_data <= "000000000000";
      when "010011010111000" => color_data <= "000000000000";
      when "010011010111001" => color_data <= "000000000000";
      when "010011010111010" => color_data <= "000000000000";
      when "010011010111011" => color_data <= "000000000000";
      when "010011010111100" => color_data <= "000000000000";
      when "010011010111101" => color_data <= "000000000000";
      when "010011010111110" => color_data <= "000000000000";
      when "010011010111111" => color_data <= "000000000000";
      when "010011011000000" => color_data <= "000000000000";
      when "010011011000001" => color_data <= "000000000000";
      when "010011011000010" => color_data <= "000000000000";
      when "010011011000011" => color_data <= "000100010001";
      when "010011011000100" => color_data <= "110010100000";
      when "010011011000101" => color_data <= "110110100000";
      when "010011011000110" => color_data <= "111110110000";
      when "010011011000111" => color_data <= "110110100000";
      when "010011011001000" => color_data <= "001000100010";
      when "010011011001001" => color_data <= "000000000000";
      when "010011011001010" => color_data <= "000000000000";
      when "010011011001011" => color_data <= "000000000000";
      when "010011011001100" => color_data <= "000000000000";
      when "010011011001101" => color_data <= "000000000000";
      when "010011011001110" => color_data <= "000000000000";
      when "010011011001111" => color_data <= "000000000000";
      when "010011011010000" => color_data <= "000000000000";
      when "010011011010001" => color_data <= "000000000000";
      when "010011011010010" => color_data <= "000000000000";
      when "010011011010011" => color_data <= "000000000000";
      when "010011011010100" => color_data <= "000000000000";
      when "010011011010101" => color_data <= "000000000000";
      when "010011011010110" => color_data <= "000000000000";
      when "010011011010111" => color_data <= "000000000000";
      when "010011011011000" => color_data <= "000000000000";
      when "010011011011001" => color_data <= "000000000000";
      when "010011011011010" => color_data <= "000000000000";
      when "010011011011011" => color_data <= "000000000000";
      when "010011011011100" => color_data <= "000000000000";
      when "010011011011101" => color_data <= "000000000000";
      when "010011011011110" => color_data <= "000000000000";
      when "010011011011111" => color_data <= "000000000000";
      when "010011011100000" => color_data <= "000000000000";
      when "010011011100001" => color_data <= "000000000000";
      when "010011011100010" => color_data <= "000000000000";
      when "010011011100011" => color_data <= "000000000000";
      when "010011100000000" => color_data <= "000000000000";
      when "010011100000001" => color_data <= "000000000000";
      when "010011100000010" => color_data <= "000000000000";
      when "010011100000011" => color_data <= "000000000000";
      when "010011100000100" => color_data <= "000000000000";
      when "010011100000101" => color_data <= "000000000000";
      when "010011100000110" => color_data <= "000000000000";
      when "010011100000111" => color_data <= "000000000000";
      when "010011100001000" => color_data <= "000000000000";
      when "010011100001001" => color_data <= "000000000000";
      when "010011100001010" => color_data <= "000000000000";
      when "010011100001011" => color_data <= "000000000000";
      when "010011100001100" => color_data <= "000000000000";
      when "010011100001101" => color_data <= "000000000000";
      when "010011100001110" => color_data <= "000000000000";
      when "010011100001111" => color_data <= "000000000000";
      when "010011100010000" => color_data <= "000000000000";
      when "010011100010001" => color_data <= "000000000000";
      when "010011100010010" => color_data <= "000000000000";
      when "010011100010011" => color_data <= "000000000000";
      when "010011100010100" => color_data <= "000000000000";
      when "010011100010101" => color_data <= "000000000000";
      when "010011100010110" => color_data <= "000000000000";
      when "010011100010111" => color_data <= "000000000000";
      when "010011100011000" => color_data <= "000000000000";
      when "010011100011001" => color_data <= "000000000000";
      when "010011100011010" => color_data <= "000000000000";
      when "010011100011011" => color_data <= "000000000000";
      when "010011100011100" => color_data <= "000000000000";
      when "010011100011101" => color_data <= "000000000000";
      when "010011100011110" => color_data <= "000000000000";
      when "010011100011111" => color_data <= "000000000000";
      when "010011100100000" => color_data <= "100110000010";
      when "010011100100001" => color_data <= "110110100000";
      when "010011100100010" => color_data <= "111110110000";
      when "010011100100011" => color_data <= "110110100000";
      when "010011100100100" => color_data <= "010000110010";
      when "010011100100101" => color_data <= "000000000000";
      when "010011100100110" => color_data <= "000000000000";
      when "010011100100111" => color_data <= "000000000000";
      when "010011100101000" => color_data <= "000000000000";
      when "010011100101001" => color_data <= "000000000000";
      when "010011100101010" => color_data <= "000000000000";
      when "010011100101011" => color_data <= "000000000000";
      when "010011100101100" => color_data <= "000000000000";
      when "010011100101101" => color_data <= "000000000000";
      when "010011100101110" => color_data <= "000000000000";
      when "010011100101111" => color_data <= "000000000000";
      when "010011100110000" => color_data <= "000000000000";
      when "010011100110001" => color_data <= "000000000000";
      when "010011100110010" => color_data <= "000000000000";
      when "010011100110011" => color_data <= "000000000000";
      when "010011100110100" => color_data <= "000000000000";
      when "010011100110101" => color_data <= "000000000000";
      when "010011100110110" => color_data <= "000000000000";
      when "010011100110111" => color_data <= "000000000000";
      when "010011100111000" => color_data <= "000000000000";
      when "010011100111001" => color_data <= "000000000000";
      when "010011100111010" => color_data <= "000000000000";
      when "010011100111011" => color_data <= "000000000000";
      when "010011100111100" => color_data <= "000000000000";
      when "010011100111101" => color_data <= "000000000000";
      when "010011100111110" => color_data <= "000000000000";
      when "010011100111111" => color_data <= "000000000000";
      when "010011101000000" => color_data <= "000000000000";
      when "010011101000001" => color_data <= "000000000000";
      when "010011101000010" => color_data <= "001100110010";
      when "010011101000011" => color_data <= "110110100000";
      when "010011101000100" => color_data <= "111110110000";
      when "010011101000101" => color_data <= "110110100000";
      when "010011101000110" => color_data <= "101110010001";
      when "010011101000111" => color_data <= "000100010001";
      when "010011101001000" => color_data <= "000000000000";
      when "010011101001001" => color_data <= "000000000000";
      when "010011101001010" => color_data <= "000000000000";
      when "010011101001011" => color_data <= "000000000000";
      when "010011101001100" => color_data <= "000000000000";
      when "010011101001101" => color_data <= "000000000000";
      when "010011101001110" => color_data <= "000000000000";
      when "010011101001111" => color_data <= "000000000000";
      when "010011101010000" => color_data <= "000000000000";
      when "010011101010001" => color_data <= "000000000000";
      when "010011101010010" => color_data <= "000000000000";
      when "010011101010011" => color_data <= "000000000000";
      when "010011101010100" => color_data <= "000000000000";
      when "010011101010101" => color_data <= "000000000000";
      when "010011101010110" => color_data <= "000000000000";
      when "010011101010111" => color_data <= "000000000000";
      when "010011101011000" => color_data <= "000000000000";
      when "010011101011001" => color_data <= "000000000000";
      when "010011101011010" => color_data <= "000000000000";
      when "010011101011011" => color_data <= "000000000000";
      when "010011101011100" => color_data <= "000000000000";
      when "010011101011101" => color_data <= "000000000000";
      when "010011101011110" => color_data <= "000000000000";
      when "010011101011111" => color_data <= "000000000000";
      when "010011101100000" => color_data <= "000000000000";
      when "010011101100001" => color_data <= "000000000000";
      when "010011101100010" => color_data <= "000000000000";
      when "010011101100011" => color_data <= "000000000000";
      when "010011110000000" => color_data <= "000000000000";
      when "010011110000001" => color_data <= "000000000000";
      when "010011110000010" => color_data <= "000000000000";
      when "010011110000011" => color_data <= "000000000000";
      when "010011110000100" => color_data <= "000000000000";
      when "010011110000101" => color_data <= "000000000000";
      when "010011110000110" => color_data <= "000000000000";
      when "010011110000111" => color_data <= "000000000000";
      when "010011110001000" => color_data <= "000000000000";
      when "010011110001001" => color_data <= "000000000000";
      when "010011110001010" => color_data <= "000000000000";
      when "010011110001011" => color_data <= "000000000000";
      when "010011110001100" => color_data <= "000000000000";
      when "010011110001101" => color_data <= "000000000000";
      when "010011110001110" => color_data <= "000000000000";
      when "010011110001111" => color_data <= "000000000000";
      when "010011110010000" => color_data <= "000000000000";
      when "010011110010001" => color_data <= "000000000000";
      when "010011110010010" => color_data <= "000000000000";
      when "010011110010011" => color_data <= "000000000000";
      when "010011110010100" => color_data <= "000000000000";
      when "010011110010101" => color_data <= "000000000000";
      when "010011110010110" => color_data <= "000000000000";
      when "010011110010111" => color_data <= "000000000000";
      when "010011110011000" => color_data <= "000000000000";
      when "010011110011001" => color_data <= "000000000000";
      when "010011110011010" => color_data <= "000000000000";
      when "010011110011011" => color_data <= "000000000000";
      when "010011110011100" => color_data <= "000000000000";
      when "010011110011101" => color_data <= "000000000000";
      when "010011110011110" => color_data <= "000000000000";
      when "010011110011111" => color_data <= "000000000000";
      when "010011110100000" => color_data <= "000000000000";
      when "010011110100001" => color_data <= "011001010011";
      when "010011110100010" => color_data <= "110110100000";
      when "010011110100011" => color_data <= "111110110000";
      when "010011110100100" => color_data <= "110110100000";
      when "010011110100101" => color_data <= "011001010011";
      when "010011110100110" => color_data <= "000000000000";
      when "010011110100111" => color_data <= "000000000000";
      when "010011110101000" => color_data <= "000000000000";
      when "010011110101001" => color_data <= "000000000000";
      when "010011110101010" => color_data <= "000000000000";
      when "010011110101011" => color_data <= "000000000000";
      when "010011110101100" => color_data <= "000000000000";
      when "010011110101101" => color_data <= "000000000000";
      when "010011110101110" => color_data <= "000000000000";
      when "010011110101111" => color_data <= "000000000000";
      when "010011110110000" => color_data <= "000000000000";
      when "010011110110001" => color_data <= "000000000000";
      when "010011110110010" => color_data <= "000000000000";
      when "010011110110011" => color_data <= "000000000000";
      when "010011110110100" => color_data <= "000000000000";
      when "010011110110101" => color_data <= "000000000000";
      when "010011110110110" => color_data <= "000000000000";
      when "010011110110111" => color_data <= "000000000000";
      when "010011110111000" => color_data <= "000000000000";
      when "010011110111001" => color_data <= "000000000000";
      when "010011110111010" => color_data <= "000000000000";
      when "010011110111011" => color_data <= "000000000000";
      when "010011110111100" => color_data <= "000000000000";
      when "010011110111101" => color_data <= "000000000000";
      when "010011110111110" => color_data <= "000000000000";
      when "010011110111111" => color_data <= "000000000000";
      when "010011111000000" => color_data <= "000000000000";
      when "010011111000001" => color_data <= "011101100011";
      when "010011111000010" => color_data <= "110110100000";
      when "010011111000011" => color_data <= "111110110000";
      when "010011111000100" => color_data <= "110110100000";
      when "010011111000101" => color_data <= "100001110010";
      when "010011111000110" => color_data <= "000000000000";
      when "010011111000111" => color_data <= "000000000000";
      when "010011111001000" => color_data <= "000000000000";
      when "010011111001001" => color_data <= "000000000000";
      when "010011111001010" => color_data <= "000000000000";
      when "010011111001011" => color_data <= "000000000000";
      when "010011111001100" => color_data <= "000000000000";
      when "010011111001101" => color_data <= "000000000000";
      when "010011111001110" => color_data <= "000000000000";
      when "010011111001111" => color_data <= "000000000000";
      when "010011111010000" => color_data <= "000000000000";
      when "010011111010001" => color_data <= "000000000000";
      when "010011111010010" => color_data <= "000000000000";
      when "010011111010011" => color_data <= "000000000000";
      when "010011111010100" => color_data <= "000000000000";
      when "010011111010101" => color_data <= "000000000000";
      when "010011111010110" => color_data <= "000000000000";
      when "010011111010111" => color_data <= "000000000000";
      when "010011111011000" => color_data <= "000000000000";
      when "010011111011001" => color_data <= "000000000000";
      when "010011111011010" => color_data <= "000000000000";
      when "010011111011011" => color_data <= "000000000000";
      when "010011111011100" => color_data <= "000000000000";
      when "010011111011101" => color_data <= "000000000000";
      when "010011111011110" => color_data <= "000000000000";
      when "010011111011111" => color_data <= "000000000000";
      when "010011111100000" => color_data <= "000000000000";
      when "010011111100001" => color_data <= "000000000000";
      when "010011111100010" => color_data <= "000000000000";
      when "010011111100011" => color_data <= "000000000000";
      when "010100000000000" => color_data <= "000000000000";
      when "010100000000001" => color_data <= "000000000000";
      when "010100000000010" => color_data <= "000000000000";
      when "010100000000011" => color_data <= "000000000000";
      when "010100000000100" => color_data <= "000000000000";
      when "010100000000101" => color_data <= "000000000000";
      when "010100000000110" => color_data <= "000000000000";
      when "010100000000111" => color_data <= "000000000000";
      when "010100000001000" => color_data <= "000000000000";
      when "010100000001001" => color_data <= "000000000000";
      when "010100000001010" => color_data <= "000000000000";
      when "010100000001011" => color_data <= "000000000000";
      when "010100000001100" => color_data <= "000000000000";
      when "010100000001101" => color_data <= "000000000000";
      when "010100000001110" => color_data <= "000000000000";
      when "010100000001111" => color_data <= "000000000000";
      when "010100000010000" => color_data <= "000000000000";
      when "010100000010001" => color_data <= "000000000000";
      when "010100000010010" => color_data <= "000000000000";
      when "010100000010011" => color_data <= "000000000000";
      when "010100000010100" => color_data <= "000000000000";
      when "010100000010101" => color_data <= "000000000000";
      when "010100000010110" => color_data <= "000000000000";
      when "010100000010111" => color_data <= "000000000000";
      when "010100000011000" => color_data <= "000000000000";
      when "010100000011001" => color_data <= "000000000000";
      when "010100000011010" => color_data <= "000000000000";
      when "010100000011011" => color_data <= "000000000000";
      when "010100000011100" => color_data <= "000000000000";
      when "010100000011101" => color_data <= "000000000000";
      when "010100000011110" => color_data <= "000000000000";
      when "010100000011111" => color_data <= "000000000000";
      when "010100000100000" => color_data <= "000000000000";
      when "010100000100001" => color_data <= "000000000000";
      when "010100000100010" => color_data <= "010000110010";
      when "010100000100011" => color_data <= "110010010000";
      when "010100000100100" => color_data <= "110110100000";
      when "010100000100101" => color_data <= "110110100000";
      when "010100000100110" => color_data <= "100101110010";
      when "010100000100111" => color_data <= "000000000000";
      when "010100000101000" => color_data <= "000000000000";
      when "010100000101001" => color_data <= "000000000000";
      when "010100000101010" => color_data <= "000000000000";
      when "010100000101011" => color_data <= "000000000000";
      when "010100000101100" => color_data <= "000000000000";
      when "010100000101101" => color_data <= "000000000000";
      when "010100000101110" => color_data <= "000000000000";
      when "010100000101111" => color_data <= "000000000000";
      when "010100000110000" => color_data <= "000000000000";
      when "010100000110001" => color_data <= "000000000000";
      when "010100000110010" => color_data <= "000000000000";
      when "010100000110011" => color_data <= "000000000000";
      when "010100000110100" => color_data <= "000000000000";
      when "010100000110101" => color_data <= "000000000000";
      when "010100000110110" => color_data <= "000000000000";
      when "010100000110111" => color_data <= "000000000000";
      when "010100000111000" => color_data <= "000000000000";
      when "010100000111001" => color_data <= "000000000000";
      when "010100000111010" => color_data <= "000000000000";
      when "010100000111011" => color_data <= "000000000000";
      when "010100000111100" => color_data <= "000000000000";
      when "010100000111101" => color_data <= "000000000000";
      when "010100000111110" => color_data <= "000000000000";
      when "010100000111111" => color_data <= "000000000000";
      when "010100001000000" => color_data <= "100110000010";
      when "010100001000001" => color_data <= "110110100000";
      when "010100001000010" => color_data <= "111110110000";
      when "010100001000011" => color_data <= "110110100000";
      when "010100001000100" => color_data <= "010101010011";
      when "010100001000101" => color_data <= "000000000000";
      when "010100001000110" => color_data <= "000000000000";
      when "010100001000111" => color_data <= "000000000000";
      when "010100001001000" => color_data <= "000000000000";
      when "010100001001001" => color_data <= "000000000000";
      when "010100001001010" => color_data <= "000000000000";
      when "010100001001011" => color_data <= "000000000000";
      when "010100001001100" => color_data <= "000000000000";
      when "010100001001101" => color_data <= "000000000000";
      when "010100001001110" => color_data <= "000000000000";
      when "010100001001111" => color_data <= "000000000000";
      when "010100001010000" => color_data <= "000000000000";
      when "010100001010001" => color_data <= "000000000000";
      when "010100001010010" => color_data <= "000000000000";
      when "010100001010011" => color_data <= "000000000000";
      when "010100001010100" => color_data <= "000000000000";
      when "010100001010101" => color_data <= "000000000000";
      when "010100001010110" => color_data <= "000000000000";
      when "010100001010111" => color_data <= "000000000000";
      when "010100001011000" => color_data <= "000000000000";
      when "010100001011001" => color_data <= "000000000000";
      when "010100001011010" => color_data <= "000000000000";
      when "010100001011011" => color_data <= "000000000000";
      when "010100001011100" => color_data <= "000000000000";
      when "010100001011101" => color_data <= "000000000000";
      when "010100001011110" => color_data <= "000000000000";
      when "010100001011111" => color_data <= "000000000000";
      when "010100001100000" => color_data <= "000000000000";
      when "010100001100001" => color_data <= "000000000000";
      when "010100001100010" => color_data <= "000000000000";
      when "010100001100011" => color_data <= "000000000000";
      when "010100010000000" => color_data <= "000000000000";
      when "010100010000001" => color_data <= "000000000000";
      when "010100010000010" => color_data <= "000000000000";
      when "010100010000011" => color_data <= "000000000000";
      when "010100010000100" => color_data <= "000000000000";
      when "010100010000101" => color_data <= "000000000000";
      when "010100010000110" => color_data <= "000000000000";
      when "010100010000111" => color_data <= "000000000000";
      when "010100010001000" => color_data <= "000000000000";
      when "010100010001001" => color_data <= "000000000000";
      when "010100010001010" => color_data <= "000000000000";
      when "010100010001011" => color_data <= "000000000000";
      when "010100010001100" => color_data <= "000000000000";
      when "010100010001101" => color_data <= "000000000000";
      when "010100010001110" => color_data <= "000000000000";
      when "010100010001111" => color_data <= "000000000000";
      when "010100010010000" => color_data <= "000000000000";
      when "010100010010001" => color_data <= "000000000000";
      when "010100010010010" => color_data <= "000000000000";
      when "010100010010011" => color_data <= "000000000000";
      when "010100010010100" => color_data <= "000000000000";
      when "010100010010101" => color_data <= "000000000000";
      when "010100010010110" => color_data <= "000000000000";
      when "010100010010111" => color_data <= "000000000000";
      when "010100010011000" => color_data <= "000000000000";
      when "010100010011001" => color_data <= "000000000000";
      when "010100010011010" => color_data <= "000000000000";
      when "010100010011011" => color_data <= "000000000000";
      when "010100010011100" => color_data <= "000000000000";
      when "010100010011101" => color_data <= "000000000000";
      when "010100010011110" => color_data <= "000000000000";
      when "010100010011111" => color_data <= "000000000000";
      when "010100010100000" => color_data <= "000000000000";
      when "010100010100001" => color_data <= "000000000000";
      when "010100010100010" => color_data <= "000000000000";
      when "010100010100011" => color_data <= "000000000000";
      when "010100010100100" => color_data <= "100101110010";
      when "010100010100101" => color_data <= "110110100000";
      when "010100010100110" => color_data <= "110110010000";
      when "010100010100111" => color_data <= "110010010001";
      when "010100010101000" => color_data <= "001100110010";
      when "010100010101001" => color_data <= "000000000000";
      when "010100010101010" => color_data <= "000000000000";
      when "010100010101011" => color_data <= "000000000000";
      when "010100010101100" => color_data <= "000000000000";
      when "010100010101101" => color_data <= "000000000000";
      when "010100010101110" => color_data <= "000000000000";
      when "010100010101111" => color_data <= "000000000000";
      when "010100010110000" => color_data <= "000000000000";
      when "010100010110001" => color_data <= "000000000000";
      when "010100010110010" => color_data <= "000000000000";
      when "010100010110011" => color_data <= "000000000000";
      when "010100010110100" => color_data <= "000000000000";
      when "010100010110101" => color_data <= "000000000000";
      when "010100010110110" => color_data <= "000000000000";
      when "010100010110111" => color_data <= "000000000000";
      when "010100010111000" => color_data <= "000000000000";
      when "010100010111001" => color_data <= "000000000000";
      when "010100010111010" => color_data <= "000000000000";
      when "010100010111011" => color_data <= "000000000000";
      when "010100010111100" => color_data <= "000000000000";
      when "010100010111101" => color_data <= "000000000000";
      when "010100010111110" => color_data <= "010001000010";
      when "010100010111111" => color_data <= "110110100000";
      when "010100011000000" => color_data <= "111110110000";
      when "010100011000001" => color_data <= "110110100000";
      when "010100011000010" => color_data <= "101010000010";
      when "010100011000011" => color_data <= "000100010001";
      when "010100011000100" => color_data <= "000000000000";
      when "010100011000101" => color_data <= "000000000000";
      when "010100011000110" => color_data <= "000000000000";
      when "010100011000111" => color_data <= "000000000000";
      when "010100011001000" => color_data <= "000000000000";
      when "010100011001001" => color_data <= "000000000000";
      when "010100011001010" => color_data <= "000000000000";
      when "010100011001011" => color_data <= "000000000000";
      when "010100011001100" => color_data <= "000000000000";
      when "010100011001101" => color_data <= "000000000000";
      when "010100011001110" => color_data <= "000000000000";
      when "010100011001111" => color_data <= "000000000000";
      when "010100011010000" => color_data <= "000000000000";
      when "010100011010001" => color_data <= "000000000000";
      when "010100011010010" => color_data <= "000000000000";
      when "010100011010011" => color_data <= "000000000000";
      when "010100011010100" => color_data <= "000000000000";
      when "010100011010101" => color_data <= "000000000000";
      when "010100011010110" => color_data <= "000000000000";
      when "010100011010111" => color_data <= "000000000000";
      when "010100011011000" => color_data <= "000000000000";
      when "010100011011001" => color_data <= "000000000000";
      when "010100011011010" => color_data <= "000000000000";
      when "010100011011011" => color_data <= "000000000000";
      when "010100011011100" => color_data <= "000000000000";
      when "010100011011101" => color_data <= "000000000000";
      when "010100011011110" => color_data <= "000000000000";
      when "010100011011111" => color_data <= "000000000000";
      when "010100011100000" => color_data <= "000000000000";
      when "010100011100001" => color_data <= "000000000000";
      when "010100011100010" => color_data <= "000000000000";
      when "010100011100011" => color_data <= "000000000000";
      when "010100100000000" => color_data <= "000000000000";
      when "010100100000001" => color_data <= "000000000000";
      when "010100100000010" => color_data <= "000000000000";
      when "010100100000011" => color_data <= "000000000000";
      when "010100100000100" => color_data <= "000000000000";
      when "010100100000101" => color_data <= "000000000000";
      when "010100100000110" => color_data <= "000000000000";
      when "010100100000111" => color_data <= "000000000000";
      when "010100100001000" => color_data <= "000000000000";
      when "010100100001001" => color_data <= "000000000000";
      when "010100100001010" => color_data <= "000000000000";
      when "010100100001011" => color_data <= "000000000000";
      when "010100100001100" => color_data <= "000000000000";
      when "010100100001101" => color_data <= "000000000000";
      when "010100100001110" => color_data <= "000000000000";
      when "010100100001111" => color_data <= "000000000000";
      when "010100100010000" => color_data <= "000000000000";
      when "010100100010001" => color_data <= "000000000000";
      when "010100100010010" => color_data <= "000000000000";
      when "010100100010011" => color_data <= "000000000000";
      when "010100100010100" => color_data <= "000000000000";
      when "010100100010101" => color_data <= "000000000000";
      when "010100100010110" => color_data <= "000000000000";
      when "010100100010111" => color_data <= "000000000000";
      when "010100100011000" => color_data <= "000000000000";
      when "010100100011001" => color_data <= "000000000000";
      when "010100100011010" => color_data <= "000000000000";
      when "010100100011011" => color_data <= "000000000000";
      when "010100100011100" => color_data <= "000000000000";
      when "010100100011101" => color_data <= "000000000000";
      when "010100100011110" => color_data <= "000000000000";
      when "010100100011111" => color_data <= "000000000000";
      when "010100100100000" => color_data <= "000000000000";
      when "010100100100001" => color_data <= "000000000000";
      when "010100100100010" => color_data <= "000000000000";
      when "010100100100011" => color_data <= "000000000000";
      when "010100100100100" => color_data <= "000000000000";
      when "010100100100101" => color_data <= "010001000010";
      when "010100100100110" => color_data <= "110010010001";
      when "010100100100111" => color_data <= "110110010000";
      when "010100100101000" => color_data <= "110110100000";
      when "010100100101001" => color_data <= "011101100011";
      when "010100100101010" => color_data <= "000000000000";
      when "010100100101011" => color_data <= "000000000000";
      when "010100100101100" => color_data <= "000000000000";
      when "010100100101101" => color_data <= "000000000000";
      when "010100100101110" => color_data <= "000000000000";
      when "010100100101111" => color_data <= "001000100001";
      when "010100100110000" => color_data <= "011001010011";
      when "010100100110001" => color_data <= "100101110010";
      when "010100100110010" => color_data <= "101010000001";
      when "010100100110011" => color_data <= "100110000010";
      when "010100100110100" => color_data <= "011101100011";
      when "010100100110101" => color_data <= "001100110010";
      when "010100100110110" => color_data <= "000000000000";
      when "010100100110111" => color_data <= "000000000000";
      when "010100100111000" => color_data <= "000000000000";
      when "010100100111001" => color_data <= "000000000000";
      when "010100100111010" => color_data <= "000000000000";
      when "010100100111011" => color_data <= "000000000000";
      when "010100100111100" => color_data <= "000000000000";
      when "010100100111101" => color_data <= "100001110010";
      when "010100100111110" => color_data <= "110110100000";
      when "010100100111111" => color_data <= "110110010000";
      when "010100101000000" => color_data <= "110010010000";
      when "010100101000001" => color_data <= "010101010011";
      when "010100101000010" => color_data <= "000000000000";
      when "010100101000011" => color_data <= "000000000000";
      when "010100101000100" => color_data <= "000000000000";
      when "010100101000101" => color_data <= "000000000000";
      when "010100101000110" => color_data <= "000000000000";
      when "010100101000111" => color_data <= "000000000000";
      when "010100101001000" => color_data <= "000000000000";
      when "010100101001001" => color_data <= "000000000000";
      when "010100101001010" => color_data <= "000000000000";
      when "010100101001011" => color_data <= "000000000000";
      when "010100101001100" => color_data <= "000000000000";
      when "010100101001101" => color_data <= "000000000000";
      when "010100101001110" => color_data <= "000000000000";
      when "010100101001111" => color_data <= "000000000000";
      when "010100101010000" => color_data <= "000000000000";
      when "010100101010001" => color_data <= "000000000000";
      when "010100101010010" => color_data <= "000000000000";
      when "010100101010011" => color_data <= "000000000000";
      when "010100101010100" => color_data <= "000000000000";
      when "010100101010101" => color_data <= "000000000000";
      when "010100101010110" => color_data <= "000000000000";
      when "010100101010111" => color_data <= "000000000000";
      when "010100101011000" => color_data <= "000000000000";
      when "010100101011001" => color_data <= "000000000000";
      when "010100101011010" => color_data <= "000000000000";
      when "010100101011011" => color_data <= "000000000000";
      when "010100101011100" => color_data <= "000000000000";
      when "010100101011101" => color_data <= "000000000000";
      when "010100101011110" => color_data <= "000000000000";
      when "010100101011111" => color_data <= "000000000000";
      when "010100101100000" => color_data <= "000000000000";
      when "010100101100001" => color_data <= "000000000000";
      when "010100101100010" => color_data <= "000000000000";
      when "010100101100011" => color_data <= "000000000000";
      when "010100110000000" => color_data <= "000000000000";
      when "010100110000001" => color_data <= "000000000000";
      when "010100110000010" => color_data <= "000000000000";
      when "010100110000011" => color_data <= "000000000000";
      when "010100110000100" => color_data <= "000000000000";
      when "010100110000101" => color_data <= "000000000000";
      when "010100110000110" => color_data <= "000000000000";
      when "010100110000111" => color_data <= "000000000000";
      when "010100110001000" => color_data <= "000000000000";
      when "010100110001001" => color_data <= "000000000000";
      when "010100110001010" => color_data <= "000000000000";
      when "010100110001011" => color_data <= "000000000000";
      when "010100110001100" => color_data <= "000000000000";
      when "010100110001101" => color_data <= "000000000000";
      when "010100110001110" => color_data <= "000000000000";
      when "010100110001111" => color_data <= "000000000000";
      when "010100110010000" => color_data <= "000000000000";
      when "010100110010001" => color_data <= "000000000000";
      when "010100110010010" => color_data <= "000000000000";
      when "010100110010011" => color_data <= "000000000000";
      when "010100110010100" => color_data <= "000000000000";
      when "010100110010101" => color_data <= "000000000000";
      when "010100110010110" => color_data <= "000000000000";
      when "010100110010111" => color_data <= "000000000000";
      when "010100110011000" => color_data <= "000000000000";
      when "010100110011001" => color_data <= "000000000000";
      when "010100110011010" => color_data <= "000000000000";
      when "010100110011011" => color_data <= "000000000000";
      when "010100110011100" => color_data <= "000000000000";
      when "010100110011101" => color_data <= "000000000000";
      when "010100110011110" => color_data <= "000000000000";
      when "010100110011111" => color_data <= "000000000000";
      when "010100110100000" => color_data <= "000000000000";
      when "010100110100001" => color_data <= "000000000000";
      when "010100110100010" => color_data <= "000000000000";
      when "010100110100011" => color_data <= "000000000000";
      when "010100110100100" => color_data <= "000000000000";
      when "010100110100101" => color_data <= "000000000000";
      when "010100110100110" => color_data <= "000000000000";
      when "010100110100111" => color_data <= "011001010011";
      when "010100110101000" => color_data <= "110110100000";
      when "010100110101001" => color_data <= "101110000000";
      when "010100110101010" => color_data <= "110110100000";
      when "010100110101011" => color_data <= "011001010011";
      when "010100110101100" => color_data <= "000000000000";
      when "010100110101101" => color_data <= "000000000000";
      when "010100110101110" => color_data <= "100110000010";
      when "010100110101111" => color_data <= "110110100000";
      when "010100110110000" => color_data <= "111110110000";
      when "010100110110001" => color_data <= "111110110000";
      when "010100110110010" => color_data <= "111111000000";
      when "010100110110011" => color_data <= "111110110000";
      when "010100110110100" => color_data <= "111110110000";
      when "010100110110101" => color_data <= "110110100000";
      when "010100110110110" => color_data <= "101110010001";
      when "010100110110111" => color_data <= "001000100001";
      when "010100110111000" => color_data <= "000000000000";
      when "010100110111001" => color_data <= "000000000000";
      when "010100110111010" => color_data <= "000000000000";
      when "010100110111011" => color_data <= "011101100011";
      when "010100110111100" => color_data <= "110110100000";
      when "010100110111101" => color_data <= "111110110000";
      when "010100110111110" => color_data <= "110110100000";
      when "010100110111111" => color_data <= "011101100011";
      when "010100111000000" => color_data <= "000000000000";
      when "010100111000001" => color_data <= "000000000000";
      when "010100111000010" => color_data <= "000000000000";
      when "010100111000011" => color_data <= "000000000000";
      when "010100111000100" => color_data <= "000000000000";
      when "010100111000101" => color_data <= "000000000000";
      when "010100111000110" => color_data <= "000000000000";
      when "010100111000111" => color_data <= "000000000000";
      when "010100111001000" => color_data <= "000000000000";
      when "010100111001001" => color_data <= "000000000000";
      when "010100111001010" => color_data <= "000000000000";
      when "010100111001011" => color_data <= "000000000000";
      when "010100111001100" => color_data <= "000000000000";
      when "010100111001101" => color_data <= "000000000000";
      when "010100111001110" => color_data <= "000000000000";
      when "010100111001111" => color_data <= "000000000000";
      when "010100111010000" => color_data <= "000000000000";
      when "010100111010001" => color_data <= "000000000000";
      when "010100111010010" => color_data <= "000000000000";
      when "010100111010011" => color_data <= "000000000000";
      when "010100111010100" => color_data <= "000000000000";
      when "010100111010101" => color_data <= "000000000000";
      when "010100111010110" => color_data <= "000000000000";
      when "010100111010111" => color_data <= "000000000000";
      when "010100111011000" => color_data <= "000000000000";
      when "010100111011001" => color_data <= "000000000000";
      when "010100111011010" => color_data <= "000000000000";
      when "010100111011011" => color_data <= "000000000000";
      when "010100111011100" => color_data <= "000000000000";
      when "010100111011101" => color_data <= "000000000000";
      when "010100111011110" => color_data <= "000000000000";
      when "010100111011111" => color_data <= "000000000000";
      when "010100111100000" => color_data <= "000000000000";
      when "010100111100001" => color_data <= "000000000000";
      when "010100111100010" => color_data <= "000000000000";
      when "010100111100011" => color_data <= "000000000000";
      when "010101000000000" => color_data <= "000000000000";
      when "010101000000001" => color_data <= "000000000000";
      when "010101000000010" => color_data <= "000000000000";
      when "010101000000011" => color_data <= "000000000000";
      when "010101000000100" => color_data <= "000000000000";
      when "010101000000101" => color_data <= "000000000000";
      when "010101000000110" => color_data <= "000000000000";
      when "010101000000111" => color_data <= "000000000000";
      when "010101000001000" => color_data <= "000000000000";
      when "010101000001001" => color_data <= "000000000000";
      when "010101000001010" => color_data <= "000000000000";
      when "010101000001011" => color_data <= "000000000000";
      when "010101000001100" => color_data <= "000000000000";
      when "010101000001101" => color_data <= "000000000000";
      when "010101000001110" => color_data <= "000000000000";
      when "010101000001111" => color_data <= "000000000000";
      when "010101000010000" => color_data <= "000000000000";
      when "010101000010001" => color_data <= "000000000000";
      when "010101000010010" => color_data <= "000000000000";
      when "010101000010011" => color_data <= "000000000000";
      when "010101000010100" => color_data <= "000000000000";
      when "010101000010101" => color_data <= "000000000000";
      when "010101000010110" => color_data <= "000000000000";
      when "010101000010111" => color_data <= "000000000000";
      when "010101000011000" => color_data <= "000000000000";
      when "010101000011001" => color_data <= "000000000000";
      when "010101000011010" => color_data <= "000000000000";
      when "010101000011011" => color_data <= "000000000000";
      when "010101000011100" => color_data <= "000000000000";
      when "010101000011101" => color_data <= "000000000000";
      when "010101000011110" => color_data <= "000000000000";
      when "010101000011111" => color_data <= "000000000000";
      when "010101000100000" => color_data <= "000000000000";
      when "010101000100001" => color_data <= "000000000000";
      when "010101000100010" => color_data <= "000000000000";
      when "010101000100011" => color_data <= "000000000000";
      when "010101000100100" => color_data <= "000000000000";
      when "010101000100101" => color_data <= "000000000000";
      when "010101000100110" => color_data <= "000000000000";
      when "010101000100111" => color_data <= "000000000000";
      when "010101000101000" => color_data <= "000000000000";
      when "010101000101001" => color_data <= "010101010011";
      when "010101000101010" => color_data <= "101010000001";
      when "010101000101011" => color_data <= "101110000000";
      when "010101000101100" => color_data <= "101010000010";
      when "010101000101101" => color_data <= "101110010001";
      when "010101000101110" => color_data <= "110110100000";
      when "010101000101111" => color_data <= "111111000001";
      when "010101000110000" => color_data <= "111111000001";
      when "010101000110001" => color_data <= "111111000001";
      when "010101000110010" => color_data <= "111111000001";
      when "010101000110011" => color_data <= "111111000001";
      when "010101000110100" => color_data <= "111111000001";
      when "010101000110101" => color_data <= "111111000001";
      when "010101000110110" => color_data <= "111110110000";
      when "010101000110111" => color_data <= "110110100000";
      when "010101000111000" => color_data <= "001100110010";
      when "010101000111001" => color_data <= "011001010011";
      when "010101000111010" => color_data <= "110110100000";
      when "010101000111011" => color_data <= "101110000000";
      when "010101000111100" => color_data <= "110010010000";
      when "010101000111101" => color_data <= "011001100011";
      when "010101000111110" => color_data <= "000000000000";
      when "010101000111111" => color_data <= "000000000000";
      when "010101001000000" => color_data <= "000000000000";
      when "010101001000001" => color_data <= "000000000000";
      when "010101001000010" => color_data <= "000000000000";
      when "010101001000011" => color_data <= "000000000000";
      when "010101001000100" => color_data <= "000000000000";
      when "010101001000101" => color_data <= "000000000000";
      when "010101001000110" => color_data <= "000000000000";
      when "010101001000111" => color_data <= "000000000000";
      when "010101001001000" => color_data <= "000000000000";
      when "010101001001001" => color_data <= "000000000000";
      when "010101001001010" => color_data <= "000000000000";
      when "010101001001011" => color_data <= "000000000000";
      when "010101001001100" => color_data <= "000000000000";
      when "010101001001101" => color_data <= "000000000000";
      when "010101001001110" => color_data <= "000000000000";
      when "010101001001111" => color_data <= "000000000000";
      when "010101001010000" => color_data <= "000000000000";
      when "010101001010001" => color_data <= "000000000000";
      when "010101001010010" => color_data <= "000000000000";
      when "010101001010011" => color_data <= "000000000000";
      when "010101001010100" => color_data <= "000000000000";
      when "010101001010101" => color_data <= "000000000000";
      when "010101001010110" => color_data <= "000000000000";
      when "010101001010111" => color_data <= "000000000000";
      when "010101001011000" => color_data <= "000000000000";
      when "010101001011001" => color_data <= "000000000000";
      when "010101001011010" => color_data <= "000000000000";
      when "010101001011011" => color_data <= "000000000000";
      when "010101001011100" => color_data <= "000000000000";
      when "010101001011101" => color_data <= "000000000000";
      when "010101001011110" => color_data <= "000000000000";
      when "010101001011111" => color_data <= "000000000000";
      when "010101001100000" => color_data <= "000000000000";
      when "010101001100001" => color_data <= "000000000000";
      when "010101001100010" => color_data <= "000000000000";
      when "010101001100011" => color_data <= "000000000000";
      when "010101010000000" => color_data <= "000000000000";
      when "010101010000001" => color_data <= "000000000000";
      when "010101010000010" => color_data <= "000000000000";
      when "010101010000011" => color_data <= "000000000000";
      when "010101010000100" => color_data <= "000000000000";
      when "010101010000101" => color_data <= "000000000000";
      when "010101010000110" => color_data <= "000000000000";
      when "010101010000111" => color_data <= "000000000000";
      when "010101010001000" => color_data <= "000000000000";
      when "010101010001001" => color_data <= "000000000000";
      when "010101010001010" => color_data <= "000000000000";
      when "010101010001011" => color_data <= "000000000000";
      when "010101010001100" => color_data <= "000000000000";
      when "010101010001101" => color_data <= "000000000000";
      when "010101010001110" => color_data <= "000000000000";
      when "010101010001111" => color_data <= "000000000000";
      when "010101010010000" => color_data <= "000000000000";
      when "010101010010001" => color_data <= "000000000000";
      when "010101010010010" => color_data <= "000000000000";
      when "010101010010011" => color_data <= "000000000000";
      when "010101010010100" => color_data <= "000000000000";
      when "010101010010101" => color_data <= "000000000000";
      when "010101010010110" => color_data <= "000000000000";
      when "010101010010111" => color_data <= "000000000000";
      when "010101010011000" => color_data <= "000000000000";
      when "010101010011001" => color_data <= "000000000000";
      when "010101010011010" => color_data <= "000000000000";
      when "010101010011011" => color_data <= "000000000000";
      when "010101010011100" => color_data <= "000000000000";
      when "010101010011101" => color_data <= "000000000000";
      when "010101010011110" => color_data <= "000000000000";
      when "010101010011111" => color_data <= "000000000000";
      when "010101010100000" => color_data <= "000000000000";
      when "010101010100001" => color_data <= "000000000000";
      when "010101010100010" => color_data <= "000000000000";
      when "010101010100011" => color_data <= "000000000000";
      when "010101010100100" => color_data <= "000000000000";
      when "010101010100101" => color_data <= "000000000000";
      when "010101010100110" => color_data <= "000000000000";
      when "010101010100111" => color_data <= "000000000000";
      when "010101010101000" => color_data <= "000000000000";
      when "010101010101001" => color_data <= "000000000000";
      when "010101010101010" => color_data <= "000000000000";
      when "010101010101011" => color_data <= "000000000000";
      when "010101010101100" => color_data <= "111111000001";
      when "010101010101101" => color_data <= "111110110000";
      when "010101010101110" => color_data <= "111111000001";
      when "010101010101111" => color_data <= "111111000001";
      when "010101010110000" => color_data <= "111111000001";
      when "010101010110001" => color_data <= "111111000001";
      when "010101010110010" => color_data <= "111111000001";
      when "010101010110011" => color_data <= "111111000001";
      when "010101010110100" => color_data <= "111111000001";
      when "010101010110101" => color_data <= "111111000001";
      when "010101010110110" => color_data <= "111111000001";
      when "010101010110111" => color_data <= "111111000000";
      when "010101010111000" => color_data <= "111110110000";
      when "010101010111001" => color_data <= "101110010001";
      when "010101010111010" => color_data <= "011001100011";
      when "010101010111011" => color_data <= "001000100001";
      when "010101010111100" => color_data <= "000000000000";
      when "010101010111101" => color_data <= "000000000000";
      when "010101010111110" => color_data <= "000000000000";
      when "010101010111111" => color_data <= "000000000000";
      when "010101011000000" => color_data <= "000000000000";
      when "010101011000001" => color_data <= "000000000000";
      when "010101011000010" => color_data <= "000000000000";
      when "010101011000011" => color_data <= "000000000000";
      when "010101011000100" => color_data <= "000000000000";
      when "010101011000101" => color_data <= "000000000000";
      when "010101011000110" => color_data <= "000000000000";
      when "010101011000111" => color_data <= "000000000000";
      when "010101011001000" => color_data <= "000000000000";
      when "010101011001001" => color_data <= "000000000000";
      when "010101011001010" => color_data <= "000000000000";
      when "010101011001011" => color_data <= "000000000000";
      when "010101011001100" => color_data <= "000000000000";
      when "010101011001101" => color_data <= "000000000000";
      when "010101011001110" => color_data <= "000000000000";
      when "010101011001111" => color_data <= "000000000000";
      when "010101011010000" => color_data <= "000000000000";
      when "010101011010001" => color_data <= "000000000000";
      when "010101011010010" => color_data <= "000000000000";
      when "010101011010011" => color_data <= "000000000000";
      when "010101011010100" => color_data <= "000000000000";
      when "010101011010101" => color_data <= "000000000000";
      when "010101011010110" => color_data <= "000000000000";
      when "010101011010111" => color_data <= "000000000000";
      when "010101011011000" => color_data <= "000000000000";
      when "010101011011001" => color_data <= "000000000000";
      when "010101011011010" => color_data <= "000000000000";
      when "010101011011011" => color_data <= "000000000000";
      when "010101011011100" => color_data <= "000000000000";
      when "010101011011101" => color_data <= "000000000000";
      when "010101011011110" => color_data <= "000000000000";
      when "010101011011111" => color_data <= "000000000000";
      when "010101011100000" => color_data <= "000000000000";
      when "010101011100001" => color_data <= "000000000000";
      when "010101011100010" => color_data <= "000000000000";
      when "010101011100011" => color_data <= "000000000000";
      when "010101100000000" => color_data <= "000000000000";
      when "010101100000001" => color_data <= "000000000000";
      when "010101100000010" => color_data <= "000000000000";
      when "010101100000011" => color_data <= "000000000000";
      when "010101100000100" => color_data <= "000000000000";
      when "010101100000101" => color_data <= "000000000000";
      when "010101100000110" => color_data <= "000000000000";
      when "010101100000111" => color_data <= "000000000000";
      when "010101100001000" => color_data <= "000000000000";
      when "010101100001001" => color_data <= "000000000000";
      when "010101100001010" => color_data <= "000000000000";
      when "010101100001011" => color_data <= "000000000000";
      when "010101100001100" => color_data <= "000000000000";
      when "010101100001101" => color_data <= "000000000000";
      when "010101100001110" => color_data <= "000000000000";
      when "010101100001111" => color_data <= "000000000000";
      when "010101100010000" => color_data <= "000000000000";
      when "010101100010001" => color_data <= "000000000000";
      when "010101100010010" => color_data <= "000000000000";
      when "010101100010011" => color_data <= "000000000000";
      when "010101100010100" => color_data <= "000000000000";
      when "010101100010101" => color_data <= "000000000000";
      when "010101100010110" => color_data <= "000000000000";
      when "010101100010111" => color_data <= "000000000000";
      when "010101100011000" => color_data <= "000000000000";
      when "010101100011001" => color_data <= "000000000000";
      when "010101100011010" => color_data <= "000000000000";
      when "010101100011011" => color_data <= "000000000000";
      when "010101100011100" => color_data <= "000000000000";
      when "010101100011101" => color_data <= "000000000000";
      when "010101100011110" => color_data <= "000000000000";
      when "010101100011111" => color_data <= "000000000000";
      when "010101100100000" => color_data <= "000000000000";
      when "010101100100001" => color_data <= "000000000000";
      when "010101100100010" => color_data <= "000000000000";
      when "010101100100011" => color_data <= "000000000000";
      when "010101100100100" => color_data <= "000000000000";
      when "010101100100101" => color_data <= "000000000000";
      when "010101100100110" => color_data <= "000000000000";
      when "010101100100111" => color_data <= "000000000000";
      when "010101100101000" => color_data <= "000000000000";
      when "010101100101001" => color_data <= "000000000000";
      when "010101100101010" => color_data <= "000000000000";
      when "010101100101011" => color_data <= "000000000000";
      when "010101100101100" => color_data <= "111111000000";
      when "010101100101101" => color_data <= "111111000000";
      when "010101100101110" => color_data <= "111111000001";
      when "010101100101111" => color_data <= "111111000001";
      when "010101100110000" => color_data <= "111111000001";
      when "010101100110001" => color_data <= "111111000001";
      when "010101100110010" => color_data <= "111111000001";
      when "010101100110011" => color_data <= "111111000001";
      when "010101100110100" => color_data <= "111111000001";
      when "010101100110101" => color_data <= "111111000001";
      when "010101100110110" => color_data <= "111111000001";
      when "010101100110111" => color_data <= "111111000001";
      when "010101100111000" => color_data <= "111110110000";
      when "010101100111001" => color_data <= "001100110010";
      when "010101100111010" => color_data <= "000000000000";
      when "010101100111011" => color_data <= "000000000000";
      when "010101100111100" => color_data <= "000000000000";
      when "010101100111101" => color_data <= "000000000000";
      when "010101100111110" => color_data <= "000000000000";
      when "010101100111111" => color_data <= "000000000000";
      when "010101101000000" => color_data <= "000000000000";
      when "010101101000001" => color_data <= "000000000000";
      when "010101101000010" => color_data <= "000000000000";
      when "010101101000011" => color_data <= "000000000000";
      when "010101101000100" => color_data <= "000000000000";
      when "010101101000101" => color_data <= "000000000000";
      when "010101101000110" => color_data <= "000000000000";
      when "010101101000111" => color_data <= "000000000000";
      when "010101101001000" => color_data <= "000000000000";
      when "010101101001001" => color_data <= "000000000000";
      when "010101101001010" => color_data <= "000000000000";
      when "010101101001011" => color_data <= "000000000000";
      when "010101101001100" => color_data <= "000000000000";
      when "010101101001101" => color_data <= "000000000000";
      when "010101101001110" => color_data <= "000000000000";
      when "010101101001111" => color_data <= "000000000000";
      when "010101101010000" => color_data <= "000000000000";
      when "010101101010001" => color_data <= "000000000000";
      when "010101101010010" => color_data <= "000000000000";
      when "010101101010011" => color_data <= "000000000000";
      when "010101101010100" => color_data <= "000000000000";
      when "010101101010101" => color_data <= "000000000000";
      when "010101101010110" => color_data <= "000000000000";
      when "010101101010111" => color_data <= "000000000000";
      when "010101101011000" => color_data <= "000000000000";
      when "010101101011001" => color_data <= "000000000000";
      when "010101101011010" => color_data <= "000000000000";
      when "010101101011011" => color_data <= "000000000000";
      when "010101101011100" => color_data <= "000000000000";
      when "010101101011101" => color_data <= "000000000000";
      when "010101101011110" => color_data <= "000000000000";
      when "010101101011111" => color_data <= "000000000000";
      when "010101101100000" => color_data <= "000000000000";
      when "010101101100001" => color_data <= "000000000000";
      when "010101101100010" => color_data <= "000000000000";
      when "010101101100011" => color_data <= "000000000000";
      when "010101110000000" => color_data <= "000000000000";
      when "010101110000001" => color_data <= "000000000000";
      when "010101110000010" => color_data <= "000000000000";
      when "010101110000011" => color_data <= "000000000000";
      when "010101110000100" => color_data <= "000000000000";
      when "010101110000101" => color_data <= "000000000000";
      when "010101110000110" => color_data <= "000000000000";
      when "010101110000111" => color_data <= "000000000000";
      when "010101110001000" => color_data <= "000000000000";
      when "010101110001001" => color_data <= "000000000000";
      when "010101110001010" => color_data <= "000000000000";
      when "010101110001011" => color_data <= "000000000000";
      when "010101110001100" => color_data <= "000000000000";
      when "010101110001101" => color_data <= "000000000000";
      when "010101110001110" => color_data <= "000000000000";
      when "010101110001111" => color_data <= "000000000000";
      when "010101110010000" => color_data <= "000000000000";
      when "010101110010001" => color_data <= "000000000000";
      when "010101110010010" => color_data <= "000000000000";
      when "010101110010011" => color_data <= "000000000000";
      when "010101110010100" => color_data <= "000000000000";
      when "010101110010101" => color_data <= "000000000000";
      when "010101110010110" => color_data <= "000000000000";
      when "010101110010111" => color_data <= "000000000000";
      when "010101110011000" => color_data <= "000000000000";
      when "010101110011001" => color_data <= "000000000000";
      when "010101110011010" => color_data <= "000000000000";
      when "010101110011011" => color_data <= "000000000000";
      when "010101110011100" => color_data <= "000000000000";
      when "010101110011101" => color_data <= "000000000000";
      when "010101110011110" => color_data <= "000000000000";
      when "010101110011111" => color_data <= "000000000000";
      when "010101110100000" => color_data <= "000000000000";
      when "010101110100001" => color_data <= "000000000000";
      when "010101110100010" => color_data <= "000000000000";
      when "010101110100011" => color_data <= "000000000000";
      when "010101110100100" => color_data <= "000000000000";
      when "010101110100101" => color_data <= "000000000000";
      when "010101110100110" => color_data <= "000000000000";
      when "010101110100111" => color_data <= "000000000000";
      when "010101110101000" => color_data <= "000000000000";
      when "010101110101001" => color_data <= "000000000000";
      when "010101110101010" => color_data <= "000000000000";
      when "010101110101011" => color_data <= "010101000010";
      when "010101110101100" => color_data <= "111110110000";
      when "010101110101101" => color_data <= "111111000001";
      when "010101110101110" => color_data <= "111111000001";
      when "010101110101111" => color_data <= "111111000001";
      when "010101110110000" => color_data <= "111111000001";
      when "010101110110001" => color_data <= "111111000001";
      when "010101110110010" => color_data <= "111111000001";
      when "010101110110011" => color_data <= "111111000001";
      when "010101110110100" => color_data <= "111111000001";
      when "010101110110101" => color_data <= "111111000001";
      when "010101110110110" => color_data <= "111111000001";
      when "010101110110111" => color_data <= "111111000001";
      when "010101110111000" => color_data <= "111110110000";
      when "010101110111001" => color_data <= "100001110010";
      when "010101110111010" => color_data <= "000000000000";
      when "010101110111011" => color_data <= "000000000000";
      when "010101110111100" => color_data <= "000000000000";
      when "010101110111101" => color_data <= "000000000000";
      when "010101110111110" => color_data <= "000000000000";
      when "010101110111111" => color_data <= "000000000000";
      when "010101111000000" => color_data <= "000000000000";
      when "010101111000001" => color_data <= "000000000000";
      when "010101111000010" => color_data <= "000000000000";
      when "010101111000011" => color_data <= "000000000000";
      when "010101111000100" => color_data <= "000000000000";
      when "010101111000101" => color_data <= "000000000000";
      when "010101111000110" => color_data <= "000000000000";
      when "010101111000111" => color_data <= "000000000000";
      when "010101111001000" => color_data <= "000000000000";
      when "010101111001001" => color_data <= "000000000000";
      when "010101111001010" => color_data <= "000000000000";
      when "010101111001011" => color_data <= "000000000000";
      when "010101111001100" => color_data <= "000000000000";
      when "010101111001101" => color_data <= "000000000000";
      when "010101111001110" => color_data <= "000000000000";
      when "010101111001111" => color_data <= "000000000000";
      when "010101111010000" => color_data <= "000000000000";
      when "010101111010001" => color_data <= "000000000000";
      when "010101111010010" => color_data <= "000000000000";
      when "010101111010011" => color_data <= "000000000000";
      when "010101111010100" => color_data <= "000000000000";
      when "010101111010101" => color_data <= "000000000000";
      when "010101111010110" => color_data <= "000000000000";
      when "010101111010111" => color_data <= "000000000000";
      when "010101111011000" => color_data <= "000000000000";
      when "010101111011001" => color_data <= "000000000000";
      when "010101111011010" => color_data <= "000000000000";
      when "010101111011011" => color_data <= "000000000000";
      when "010101111011100" => color_data <= "000000000000";
      when "010101111011101" => color_data <= "000000000000";
      when "010101111011110" => color_data <= "000000000000";
      when "010101111011111" => color_data <= "000000000000";
      when "010101111100000" => color_data <= "000000000000";
      when "010101111100001" => color_data <= "000000000000";
      when "010101111100010" => color_data <= "000000000000";
      when "010101111100011" => color_data <= "000000000000";
      when "010110000000000" => color_data <= "000000000000";
      when "010110000000001" => color_data <= "000000000000";
      when "010110000000010" => color_data <= "000000000000";
      when "010110000000011" => color_data <= "000000000000";
      when "010110000000100" => color_data <= "000000000000";
      when "010110000000101" => color_data <= "000000000000";
      when "010110000000110" => color_data <= "000000000000";
      when "010110000000111" => color_data <= "000000000000";
      when "010110000001000" => color_data <= "000000000000";
      when "010110000001001" => color_data <= "000000000000";
      when "010110000001010" => color_data <= "000000000000";
      when "010110000001011" => color_data <= "000000000000";
      when "010110000001100" => color_data <= "000000000000";
      when "010110000001101" => color_data <= "000000000000";
      when "010110000001110" => color_data <= "000000000000";
      when "010110000001111" => color_data <= "000000000000";
      when "010110000010000" => color_data <= "000000000000";
      when "010110000010001" => color_data <= "000000000000";
      when "010110000010010" => color_data <= "000000000000";
      when "010110000010011" => color_data <= "000000000000";
      when "010110000010100" => color_data <= "000000000000";
      when "010110000010101" => color_data <= "000000000000";
      when "010110000010110" => color_data <= "000000000000";
      when "010110000010111" => color_data <= "000000000000";
      when "010110000011000" => color_data <= "000000000000";
      when "010110000011001" => color_data <= "000000000000";
      when "010110000011010" => color_data <= "000000000000";
      when "010110000011011" => color_data <= "000000000000";
      when "010110000011100" => color_data <= "000000000000";
      when "010110000011101" => color_data <= "000000000000";
      when "010110000011110" => color_data <= "000000000000";
      when "010110000011111" => color_data <= "000000000000";
      when "010110000100000" => color_data <= "000000000000";
      when "010110000100001" => color_data <= "000000000000";
      when "010110000100010" => color_data <= "000000000000";
      when "010110000100011" => color_data <= "000000000000";
      when "010110000100100" => color_data <= "000000000000";
      when "010110000100101" => color_data <= "000000000000";
      when "010110000100110" => color_data <= "000000000000";
      when "010110000100111" => color_data <= "000000000000";
      when "010110000101000" => color_data <= "000000000000";
      when "010110000101001" => color_data <= "000000000000";
      when "010110000101010" => color_data <= "000000000000";
      when "010110000101011" => color_data <= "010001000010";
      when "010110000101100" => color_data <= "111110110000";
      when "010110000101101" => color_data <= "111111000001";
      when "010110000101110" => color_data <= "111111000001";
      when "010110000101111" => color_data <= "111111000001";
      when "010110000110000" => color_data <= "111111000001";
      when "010110000110001" => color_data <= "111111000001";
      when "010110000110010" => color_data <= "111111000001";
      when "010110000110011" => color_data <= "111111000001";
      when "010110000110100" => color_data <= "111111000001";
      when "010110000110101" => color_data <= "111111000001";
      when "010110000110110" => color_data <= "111111000001";
      when "010110000110111" => color_data <= "111111000001";
      when "010110000111000" => color_data <= "111110110000";
      when "010110000111001" => color_data <= "011101100011";
      when "010110000111010" => color_data <= "000000000000";
      when "010110000111011" => color_data <= "000000000000";
      when "010110000111100" => color_data <= "000000000000";
      when "010110000111101" => color_data <= "000000000000";
      when "010110000111110" => color_data <= "000000000000";
      when "010110000111111" => color_data <= "000000000000";
      when "010110001000000" => color_data <= "000000000000";
      when "010110001000001" => color_data <= "000000000000";
      when "010110001000010" => color_data <= "000000000000";
      when "010110001000011" => color_data <= "000000000000";
      when "010110001000100" => color_data <= "000000000000";
      when "010110001000101" => color_data <= "000000000000";
      when "010110001000110" => color_data <= "000000000000";
      when "010110001000111" => color_data <= "000000000000";
      when "010110001001000" => color_data <= "000000000000";
      when "010110001001001" => color_data <= "000000000000";
      when "010110001001010" => color_data <= "000000000000";
      when "010110001001011" => color_data <= "000000000000";
      when "010110001001100" => color_data <= "000000000000";
      when "010110001001101" => color_data <= "000000000000";
      when "010110001001110" => color_data <= "000000000000";
      when "010110001001111" => color_data <= "000000000000";
      when "010110001010000" => color_data <= "000000000000";
      when "010110001010001" => color_data <= "000000000000";
      when "010110001010010" => color_data <= "000000000000";
      when "010110001010011" => color_data <= "000000000000";
      when "010110001010100" => color_data <= "000000000000";
      when "010110001010101" => color_data <= "000000000000";
      when "010110001010110" => color_data <= "000000000000";
      when "010110001010111" => color_data <= "000000000000";
      when "010110001011000" => color_data <= "000000000000";
      when "010110001011001" => color_data <= "000000000000";
      when "010110001011010" => color_data <= "000000000000";
      when "010110001011011" => color_data <= "000000000000";
      when "010110001011100" => color_data <= "000000000000";
      when "010110001011101" => color_data <= "000000000000";
      when "010110001011110" => color_data <= "000000000000";
      when "010110001011111" => color_data <= "000000000000";
      when "010110001100000" => color_data <= "000000000000";
      when "010110001100001" => color_data <= "000000000000";
      when "010110001100010" => color_data <= "000000000000";
      when "010110001100011" => color_data <= "000000000000";
      when "010110010000000" => color_data <= "000000000000";
      when "010110010000001" => color_data <= "000000000000";
      when "010110010000010" => color_data <= "000000000000";
      when "010110010000011" => color_data <= "000000000000";
      when "010110010000100" => color_data <= "000000000000";
      when "010110010000101" => color_data <= "000000000000";
      when "010110010000110" => color_data <= "000000000000";
      when "010110010000111" => color_data <= "000000000000";
      when "010110010001000" => color_data <= "000000000000";
      when "010110010001001" => color_data <= "000000000000";
      when "010110010001010" => color_data <= "000000000000";
      when "010110010001011" => color_data <= "000000000000";
      when "010110010001100" => color_data <= "000000000000";
      when "010110010001101" => color_data <= "000000000000";
      when "010110010001110" => color_data <= "000000000000";
      when "010110010001111" => color_data <= "000000000000";
      when "010110010010000" => color_data <= "000000000000";
      when "010110010010001" => color_data <= "000000000000";
      when "010110010010010" => color_data <= "000000000000";
      when "010110010010011" => color_data <= "000000000000";
      when "010110010010100" => color_data <= "000000000000";
      when "010110010010101" => color_data <= "000000000000";
      when "010110010010110" => color_data <= "000000000000";
      when "010110010010111" => color_data <= "000000000000";
      when "010110010011000" => color_data <= "000000000000";
      when "010110010011001" => color_data <= "000000000000";
      when "010110010011010" => color_data <= "000000000000";
      when "010110010011011" => color_data <= "000000000000";
      when "010110010011100" => color_data <= "000000000000";
      when "010110010011101" => color_data <= "000000000000";
      when "010110010011110" => color_data <= "000000000000";
      when "010110010011111" => color_data <= "000000000000";
      when "010110010100000" => color_data <= "000000000000";
      when "010110010100001" => color_data <= "000000000000";
      when "010110010100010" => color_data <= "000000000000";
      when "010110010100011" => color_data <= "000000000000";
      when "010110010100100" => color_data <= "000000000000";
      when "010110010100101" => color_data <= "000000000000";
      when "010110010100110" => color_data <= "000000000000";
      when "010110010100111" => color_data <= "000000000000";
      when "010110010101000" => color_data <= "000000000000";
      when "010110010101001" => color_data <= "000000000000";
      when "010110010101010" => color_data <= "000000000000";
      when "010110010101011" => color_data <= "000000000000";
      when "010110010101100" => color_data <= "110110100000";
      when "010110010101101" => color_data <= "111111000000";
      when "010110010101110" => color_data <= "111111000001";
      when "010110010101111" => color_data <= "111111000001";
      when "010110010110000" => color_data <= "111111000001";
      when "010110010110001" => color_data <= "111111000001";
      when "010110010110010" => color_data <= "111111000001";
      when "010110010110011" => color_data <= "111111000001";
      when "010110010110100" => color_data <= "111111000001";
      when "010110010110101" => color_data <= "111111000001";
      when "010110010110110" => color_data <= "111111000001";
      when "010110010110111" => color_data <= "111111000001";
      when "010110010111000" => color_data <= "110110100000";
      when "010110010111001" => color_data <= "001100110010";
      when "010110010111010" => color_data <= "000000000000";
      when "010110010111011" => color_data <= "000000000000";
      when "010110010111100" => color_data <= "000000000000";
      when "010110010111101" => color_data <= "000000000000";
      when "010110010111110" => color_data <= "000000000000";
      when "010110010111111" => color_data <= "000000000000";
      when "010110011000000" => color_data <= "000000000000";
      when "010110011000001" => color_data <= "000000000000";
      when "010110011000010" => color_data <= "000000000000";
      when "010110011000011" => color_data <= "000000000000";
      when "010110011000100" => color_data <= "000000000000";
      when "010110011000101" => color_data <= "000000000000";
      when "010110011000110" => color_data <= "000000000000";
      when "010110011000111" => color_data <= "000000000000";
      when "010110011001000" => color_data <= "000000000000";
      when "010110011001001" => color_data <= "000000000000";
      when "010110011001010" => color_data <= "000000000000";
      when "010110011001011" => color_data <= "000000000000";
      when "010110011001100" => color_data <= "000000000000";
      when "010110011001101" => color_data <= "000000000000";
      when "010110011001110" => color_data <= "000000000000";
      when "010110011001111" => color_data <= "000000000000";
      when "010110011010000" => color_data <= "000000000000";
      when "010110011010001" => color_data <= "000000000000";
      when "010110011010010" => color_data <= "000000000000";
      when "010110011010011" => color_data <= "000000000000";
      when "010110011010100" => color_data <= "000000000000";
      when "010110011010101" => color_data <= "000000000000";
      when "010110011010110" => color_data <= "000000000000";
      when "010110011010111" => color_data <= "000000000000";
      when "010110011011000" => color_data <= "000000000000";
      when "010110011011001" => color_data <= "000000000000";
      when "010110011011010" => color_data <= "000000000000";
      when "010110011011011" => color_data <= "000000000000";
      when "010110011011100" => color_data <= "000000000000";
      when "010110011011101" => color_data <= "000000000000";
      when "010110011011110" => color_data <= "000000000000";
      when "010110011011111" => color_data <= "000000000000";
      when "010110011100000" => color_data <= "000000000000";
      when "010110011100001" => color_data <= "000000000000";
      when "010110011100010" => color_data <= "000000000000";
      when "010110011100011" => color_data <= "000000000000";
      when "010110100000000" => color_data <= "000000000000";
      when "010110100000001" => color_data <= "000000000000";
      when "010110100000010" => color_data <= "000000000000";
      when "010110100000011" => color_data <= "000000000000";
      when "010110100000100" => color_data <= "000000000000";
      when "010110100000101" => color_data <= "000000000000";
      when "010110100000110" => color_data <= "000000000000";
      when "010110100000111" => color_data <= "000000000000";
      when "010110100001000" => color_data <= "000000000000";
      when "010110100001001" => color_data <= "000000000000";
      when "010110100001010" => color_data <= "000000000000";
      when "010110100001011" => color_data <= "000000000000";
      when "010110100001100" => color_data <= "000000000000";
      when "010110100001101" => color_data <= "000000000000";
      when "010110100001110" => color_data <= "000000000000";
      when "010110100001111" => color_data <= "000000000000";
      when "010110100010000" => color_data <= "000000000000";
      when "010110100010001" => color_data <= "000000000000";
      when "010110100010010" => color_data <= "000000000000";
      when "010110100010011" => color_data <= "000000000000";
      when "010110100010100" => color_data <= "000000000000";
      when "010110100010101" => color_data <= "000000000000";
      when "010110100010110" => color_data <= "000000000000";
      when "010110100010111" => color_data <= "000000000000";
      when "010110100011000" => color_data <= "000000000000";
      when "010110100011001" => color_data <= "000000000000";
      when "010110100011010" => color_data <= "000000000000";
      when "010110100011011" => color_data <= "000000000000";
      when "010110100011100" => color_data <= "000000000000";
      when "010110100011101" => color_data <= "000000000000";
      when "010110100011110" => color_data <= "000000000000";
      when "010110100011111" => color_data <= "000000000000";
      when "010110100100000" => color_data <= "000000000000";
      when "010110100100001" => color_data <= "000000000000";
      when "010110100100010" => color_data <= "000000000000";
      when "010110100100011" => color_data <= "000000000000";
      when "010110100100100" => color_data <= "000000000000";
      when "010110100100101" => color_data <= "000000000000";
      when "010110100100110" => color_data <= "000000000000";
      when "010110100100111" => color_data <= "000000000000";
      when "010110100101000" => color_data <= "000000000000";
      when "010110100101001" => color_data <= "000000000000";
      when "010110100101010" => color_data <= "000000000000";
      when "010110100101011" => color_data <= "000000000000";
      when "010110100101100" => color_data <= "011001010011";
      when "010110100101101" => color_data <= "110110010000";
      when "010110100101110" => color_data <= "111111000000";
      when "010110100101111" => color_data <= "111111000001";
      when "010110100110000" => color_data <= "111111000001";
      when "010110100110001" => color_data <= "111111000001";
      when "010110100110010" => color_data <= "111111000001";
      when "010110100110011" => color_data <= "111111000001";
      when "010110100110100" => color_data <= "111111000001";
      when "010110100110101" => color_data <= "111111000001";
      when "010110100110110" => color_data <= "111111000001";
      when "010110100110111" => color_data <= "110110100000";
      when "010110100111000" => color_data <= "101010000010";
      when "010110100111001" => color_data <= "000000000000";
      when "010110100111010" => color_data <= "000000000000";
      when "010110100111011" => color_data <= "000000000000";
      when "010110100111100" => color_data <= "000000000000";
      when "010110100111101" => color_data <= "000000000000";
      when "010110100111110" => color_data <= "000000000000";
      when "010110100111111" => color_data <= "000000000000";
      when "010110101000000" => color_data <= "000000000000";
      when "010110101000001" => color_data <= "000000000000";
      when "010110101000010" => color_data <= "000000000000";
      when "010110101000011" => color_data <= "000000000000";
      when "010110101000100" => color_data <= "000000000000";
      when "010110101000101" => color_data <= "000000000000";
      when "010110101000110" => color_data <= "000000000000";
      when "010110101000111" => color_data <= "000000000000";
      when "010110101001000" => color_data <= "000000000000";
      when "010110101001001" => color_data <= "000000000000";
      when "010110101001010" => color_data <= "000000000000";
      when "010110101001011" => color_data <= "000000000000";
      when "010110101001100" => color_data <= "000000000000";
      when "010110101001101" => color_data <= "000000000000";
      when "010110101001110" => color_data <= "000000000000";
      when "010110101001111" => color_data <= "000000000000";
      when "010110101010000" => color_data <= "000000000000";
      when "010110101010001" => color_data <= "000000000000";
      when "010110101010010" => color_data <= "000000000000";
      when "010110101010011" => color_data <= "000000000000";
      when "010110101010100" => color_data <= "000000000000";
      when "010110101010101" => color_data <= "000000000000";
      when "010110101010110" => color_data <= "000000000000";
      when "010110101010111" => color_data <= "000000000000";
      when "010110101011000" => color_data <= "000000000000";
      when "010110101011001" => color_data <= "000000000000";
      when "010110101011010" => color_data <= "000000000000";
      when "010110101011011" => color_data <= "000000000000";
      when "010110101011100" => color_data <= "000000000000";
      when "010110101011101" => color_data <= "000000000000";
      when "010110101011110" => color_data <= "000000000000";
      when "010110101011111" => color_data <= "000000000000";
      when "010110101100000" => color_data <= "000000000000";
      when "010110101100001" => color_data <= "000000000000";
      when "010110101100010" => color_data <= "000000000000";
      when "010110101100011" => color_data <= "000000000000";
      when "010110110000000" => color_data <= "000000000000";
      when "010110110000001" => color_data <= "000000000000";
      when "010110110000010" => color_data <= "000000000000";
      when "010110110000011" => color_data <= "000000000000";
      when "010110110000100" => color_data <= "000000000000";
      when "010110110000101" => color_data <= "000000000000";
      when "010110110000110" => color_data <= "000000000000";
      when "010110110000111" => color_data <= "000000000000";
      when "010110110001000" => color_data <= "000000000000";
      when "010110110001001" => color_data <= "000000000000";
      when "010110110001010" => color_data <= "000000000000";
      when "010110110001011" => color_data <= "000000000000";
      when "010110110001100" => color_data <= "000000000000";
      when "010110110001101" => color_data <= "000000000000";
      when "010110110001110" => color_data <= "000000000000";
      when "010110110001111" => color_data <= "000000000000";
      when "010110110010000" => color_data <= "000000000000";
      when "010110110010001" => color_data <= "000000000000";
      when "010110110010010" => color_data <= "000000000000";
      when "010110110010011" => color_data <= "000000000000";
      when "010110110010100" => color_data <= "000000000000";
      when "010110110010101" => color_data <= "000000000000";
      when "010110110010110" => color_data <= "000000000000";
      when "010110110010111" => color_data <= "000000000000";
      when "010110110011000" => color_data <= "000000000000";
      when "010110110011001" => color_data <= "000000000000";
      when "010110110011010" => color_data <= "000000000000";
      when "010110110011011" => color_data <= "000000000000";
      when "010110110011100" => color_data <= "000000000000";
      when "010110110011101" => color_data <= "000000000000";
      when "010110110011110" => color_data <= "000000000000";
      when "010110110011111" => color_data <= "000000000000";
      when "010110110100000" => color_data <= "000000000000";
      when "010110110100001" => color_data <= "000000000000";
      when "010110110100010" => color_data <= "000000000000";
      when "010110110100011" => color_data <= "000000000000";
      when "010110110100100" => color_data <= "000000000000";
      when "010110110100101" => color_data <= "000000000000";
      when "010110110100110" => color_data <= "000000000000";
      when "010110110100111" => color_data <= "000000000000";
      when "010110110101000" => color_data <= "000000000000";
      when "010110110101001" => color_data <= "000000000000";
      when "010110110101010" => color_data <= "000000000000";
      when "010110110101011" => color_data <= "000000000000";
      when "010110110101100" => color_data <= "000000000000";
      when "010110110101101" => color_data <= "100001110010";
      when "010110110101110" => color_data <= "110110100000";
      when "010110110101111" => color_data <= "111111000001";
      when "010110110110000" => color_data <= "111111000001";
      when "010110110110001" => color_data <= "111111000001";
      when "010110110110010" => color_data <= "111111000001";
      when "010110110110011" => color_data <= "111111000001";
      when "010110110110100" => color_data <= "111111000001";
      when "010110110110101" => color_data <= "111111000001";
      when "010110110110110" => color_data <= "110110100000";
      when "010110110110111" => color_data <= "101010000010";
      when "010110110111000" => color_data <= "000000000000";
      when "010110110111001" => color_data <= "000000000000";
      when "010110110111010" => color_data <= "000000000000";
      when "010110110111011" => color_data <= "000000000000";
      when "010110110111100" => color_data <= "000000000000";
      when "010110110111101" => color_data <= "000000000000";
      when "010110110111110" => color_data <= "000000000000";
      when "010110110111111" => color_data <= "000000000000";
      when "010110111000000" => color_data <= "000000000000";
      when "010110111000001" => color_data <= "000000000000";
      when "010110111000010" => color_data <= "000000000000";
      when "010110111000011" => color_data <= "000000000000";
      when "010110111000100" => color_data <= "000000000000";
      when "010110111000101" => color_data <= "000000000000";
      when "010110111000110" => color_data <= "000000000000";
      when "010110111000111" => color_data <= "000000000000";
      when "010110111001000" => color_data <= "000000000000";
      when "010110111001001" => color_data <= "000000000000";
      when "010110111001010" => color_data <= "000000000000";
      when "010110111001011" => color_data <= "000000000000";
      when "010110111001100" => color_data <= "000000000000";
      when "010110111001101" => color_data <= "000000000000";
      when "010110111001110" => color_data <= "000000000000";
      when "010110111001111" => color_data <= "000000000000";
      when "010110111010000" => color_data <= "000000000000";
      when "010110111010001" => color_data <= "000000000000";
      when "010110111010010" => color_data <= "000000000000";
      when "010110111010011" => color_data <= "000000000000";
      when "010110111010100" => color_data <= "000000000000";
      when "010110111010101" => color_data <= "000000000000";
      when "010110111010110" => color_data <= "000000000000";
      when "010110111010111" => color_data <= "000000000000";
      when "010110111011000" => color_data <= "000000000000";
      when "010110111011001" => color_data <= "000000000000";
      when "010110111011010" => color_data <= "000000000000";
      when "010110111011011" => color_data <= "000000000000";
      when "010110111011100" => color_data <= "000000000000";
      when "010110111011101" => color_data <= "000000000000";
      when "010110111011110" => color_data <= "000000000000";
      when "010110111011111" => color_data <= "000000000000";
      when "010110111100000" => color_data <= "000000000000";
      when "010110111100001" => color_data <= "000000000000";
      when "010110111100010" => color_data <= "000000000000";
      when "010110111100011" => color_data <= "000000000000";
      when "010111000000000" => color_data <= "000000000000";
      when "010111000000001" => color_data <= "000000000000";
      when "010111000000010" => color_data <= "000000000000";
      when "010111000000011" => color_data <= "000000000000";
      when "010111000000100" => color_data <= "000000000000";
      when "010111000000101" => color_data <= "000000000000";
      when "010111000000110" => color_data <= "000000000000";
      when "010111000000111" => color_data <= "000000000000";
      when "010111000001000" => color_data <= "000000000000";
      when "010111000001001" => color_data <= "000000000000";
      when "010111000001010" => color_data <= "000000000000";
      when "010111000001011" => color_data <= "000000000000";
      when "010111000001100" => color_data <= "000000000000";
      when "010111000001101" => color_data <= "000000000000";
      when "010111000001110" => color_data <= "000000000000";
      when "010111000001111" => color_data <= "000000000000";
      when "010111000010000" => color_data <= "000000000000";
      when "010111000010001" => color_data <= "000000000000";
      when "010111000010010" => color_data <= "000000000000";
      when "010111000010011" => color_data <= "000000000000";
      when "010111000010100" => color_data <= "000000000000";
      when "010111000010101" => color_data <= "000000000000";
      when "010111000010110" => color_data <= "000000000000";
      when "010111000010111" => color_data <= "000000000000";
      when "010111000011000" => color_data <= "000000000000";
      when "010111000011001" => color_data <= "000000000000";
      when "010111000011010" => color_data <= "000000000000";
      when "010111000011011" => color_data <= "000000000000";
      when "010111000011100" => color_data <= "000000000000";
      when "010111000011101" => color_data <= "000000000000";
      when "010111000011110" => color_data <= "000000000000";
      when "010111000011111" => color_data <= "000000000000";
      when "010111000100000" => color_data <= "000000000000";
      when "010111000100001" => color_data <= "000000000000";
      when "010111000100010" => color_data <= "000000000000";
      when "010111000100011" => color_data <= "000000000000";
      when "010111000100100" => color_data <= "000000000000";
      when "010111000100101" => color_data <= "000000000000";
      when "010111000100110" => color_data <= "000000000000";
      when "010111000100111" => color_data <= "000000000000";
      when "010111000101000" => color_data <= "000000000000";
      when "010111000101001" => color_data <= "000000000000";
      when "010111000101010" => color_data <= "000000000000";
      when "010111000101011" => color_data <= "000000000000";
      when "010111000101100" => color_data <= "000000000000";
      when "010111000101101" => color_data <= "000000000000";
      when "010111000101110" => color_data <= "011001010011";
      when "010111000101111" => color_data <= "111110110000";
      when "010111000110000" => color_data <= "111111000001";
      when "010111000110001" => color_data <= "111111000001";
      when "010111000110010" => color_data <= "111111000001";
      when "010111000110011" => color_data <= "111111000001";
      when "010111000110100" => color_data <= "111111000001";
      when "010111000110101" => color_data <= "111111000000";
      when "010111000110110" => color_data <= "101010000010";
      when "010111000110111" => color_data <= "000000000000";
      when "010111000111000" => color_data <= "000000000000";
      when "010111000111001" => color_data <= "000000000000";
      when "010111000111010" => color_data <= "000000000000";
      when "010111000111011" => color_data <= "000000000000";
      when "010111000111100" => color_data <= "000000000000";
      when "010111000111101" => color_data <= "000000000000";
      when "010111000111110" => color_data <= "000000000000";
      when "010111000111111" => color_data <= "000000000000";
      when "010111001000000" => color_data <= "000000000000";
      when "010111001000001" => color_data <= "000000000000";
      when "010111001000010" => color_data <= "000000000000";
      when "010111001000011" => color_data <= "000000000000";
      when "010111001000100" => color_data <= "000000000000";
      when "010111001000101" => color_data <= "000000000000";
      when "010111001000110" => color_data <= "000000000000";
      when "010111001000111" => color_data <= "000000000000";
      when "010111001001000" => color_data <= "000000000000";
      when "010111001001001" => color_data <= "000000000000";
      when "010111001001010" => color_data <= "000000000000";
      when "010111001001011" => color_data <= "000000000000";
      when "010111001001100" => color_data <= "000000000000";
      when "010111001001101" => color_data <= "000000000000";
      when "010111001001110" => color_data <= "000000000000";
      when "010111001001111" => color_data <= "000000000000";
      when "010111001010000" => color_data <= "000000000000";
      when "010111001010001" => color_data <= "000000000000";
      when "010111001010010" => color_data <= "000000000000";
      when "010111001010011" => color_data <= "000000000000";
      when "010111001010100" => color_data <= "000000000000";
      when "010111001010101" => color_data <= "000000000000";
      when "010111001010110" => color_data <= "000000000000";
      when "010111001010111" => color_data <= "000000000000";
      when "010111001011000" => color_data <= "000000000000";
      when "010111001011001" => color_data <= "000000000000";
      when "010111001011010" => color_data <= "000000000000";
      when "010111001011011" => color_data <= "000000000000";
      when "010111001011100" => color_data <= "000000000000";
      when "010111001011101" => color_data <= "000000000000";
      when "010111001011110" => color_data <= "000000000000";
      when "010111001011111" => color_data <= "000000000000";
      when "010111001100000" => color_data <= "000000000000";
      when "010111001100001" => color_data <= "000000000000";
      when "010111001100010" => color_data <= "000000000000";
      when "010111001100011" => color_data <= "000000000000";
      when "010111010000000" => color_data <= "000000000000";
      when "010111010000001" => color_data <= "000000000000";
      when "010111010000010" => color_data <= "000000000000";
      when "010111010000011" => color_data <= "000000000000";
      when "010111010000100" => color_data <= "000000000000";
      when "010111010000101" => color_data <= "000000000000";
      when "010111010000110" => color_data <= "000000000000";
      when "010111010000111" => color_data <= "000000000000";
      when "010111010001000" => color_data <= "000000000000";
      when "010111010001001" => color_data <= "000000000000";
      when "010111010001010" => color_data <= "000000000000";
      when "010111010001011" => color_data <= "000000000000";
      when "010111010001100" => color_data <= "000000000000";
      when "010111010001101" => color_data <= "000000000000";
      when "010111010001110" => color_data <= "000000000000";
      when "010111010001111" => color_data <= "000000000000";
      when "010111010010000" => color_data <= "000000000000";
      when "010111010010001" => color_data <= "000000000000";
      when "010111010010010" => color_data <= "000000000000";
      when "010111010010011" => color_data <= "000000000000";
      when "010111010010100" => color_data <= "000000000000";
      when "010111010010101" => color_data <= "000000000000";
      when "010111010010110" => color_data <= "000000000000";
      when "010111010010111" => color_data <= "000000000000";
      when "010111010011000" => color_data <= "000000000000";
      when "010111010011001" => color_data <= "000000000000";
      when "010111010011010" => color_data <= "000000000000";
      when "010111010011011" => color_data <= "000000000000";
      when "010111010011100" => color_data <= "000000000000";
      when "010111010011101" => color_data <= "000000000000";
      when "010111010011110" => color_data <= "000000000000";
      when "010111010011111" => color_data <= "000000000000";
      when "010111010100000" => color_data <= "000000000000";
      when "010111010100001" => color_data <= "000000000000";
      when "010111010100010" => color_data <= "000000000000";
      when "010111010100011" => color_data <= "000000000000";
      when "010111010100100" => color_data <= "000000000000";
      when "010111010100101" => color_data <= "000000000000";
      when "010111010100110" => color_data <= "000000000000";
      when "010111010100111" => color_data <= "000000000000";
      when "010111010101000" => color_data <= "000000000000";
      when "010111010101001" => color_data <= "000000000000";
      when "010111010101010" => color_data <= "000000000000";
      when "010111010101011" => color_data <= "000000000000";
      when "010111010101100" => color_data <= "000000000000";
      when "010111010101101" => color_data <= "000000000000";
      when "010111010101110" => color_data <= "000100010001";
      when "010111010101111" => color_data <= "111110110000";
      when "010111010110000" => color_data <= "111111000001";
      when "010111010110001" => color_data <= "111111000001";
      when "010111010110010" => color_data <= "111111000001";
      when "010111010110011" => color_data <= "111111000001";
      when "010111010110100" => color_data <= "111111000001";
      when "010111010110101" => color_data <= "111110110000";
      when "010111010110110" => color_data <= "011101100011";
      when "010111010110111" => color_data <= "000000000000";
      when "010111010111000" => color_data <= "000000000000";
      when "010111010111001" => color_data <= "000000000000";
      when "010111010111010" => color_data <= "000000000000";
      when "010111010111011" => color_data <= "000000000000";
      when "010111010111100" => color_data <= "000000000000";
      when "010111010111101" => color_data <= "000000000000";
      when "010111010111110" => color_data <= "000000000000";
      when "010111010111111" => color_data <= "000000000000";
      when "010111011000000" => color_data <= "000000000000";
      when "010111011000001" => color_data <= "000000000000";
      when "010111011000010" => color_data <= "000000000000";
      when "010111011000011" => color_data <= "000000000000";
      when "010111011000100" => color_data <= "000000000000";
      when "010111011000101" => color_data <= "000000000000";
      when "010111011000110" => color_data <= "000000000000";
      when "010111011000111" => color_data <= "000000000000";
      when "010111011001000" => color_data <= "000000000000";
      when "010111011001001" => color_data <= "000000000000";
      when "010111011001010" => color_data <= "000000000000";
      when "010111011001011" => color_data <= "000000000000";
      when "010111011001100" => color_data <= "000000000000";
      when "010111011001101" => color_data <= "000000000000";
      when "010111011001110" => color_data <= "000000000000";
      when "010111011001111" => color_data <= "000000000000";
      when "010111011010000" => color_data <= "000000000000";
      when "010111011010001" => color_data <= "000000000000";
      when "010111011010010" => color_data <= "000000000000";
      when "010111011010011" => color_data <= "000000000000";
      when "010111011010100" => color_data <= "000000000000";
      when "010111011010101" => color_data <= "000000000000";
      when "010111011010110" => color_data <= "000000000000";
      when "010111011010111" => color_data <= "000000000000";
      when "010111011011000" => color_data <= "000000000000";
      when "010111011011001" => color_data <= "000000000000";
      when "010111011011010" => color_data <= "000000000000";
      when "010111011011011" => color_data <= "000000000000";
      when "010111011011100" => color_data <= "000000000000";
      when "010111011011101" => color_data <= "000000000000";
      when "010111011011110" => color_data <= "000000000000";
      when "010111011011111" => color_data <= "000000000000";
      when "010111011100000" => color_data <= "000000000000";
      when "010111011100001" => color_data <= "000000000000";
      when "010111011100010" => color_data <= "000000000000";
      when "010111011100011" => color_data <= "000000000000";
      when "010111100000000" => color_data <= "000000000000";
      when "010111100000001" => color_data <= "000000000000";
      when "010111100000010" => color_data <= "000000000000";
      when "010111100000011" => color_data <= "000000000000";
      when "010111100000100" => color_data <= "000000000000";
      when "010111100000101" => color_data <= "000000000000";
      when "010111100000110" => color_data <= "000000000000";
      when "010111100000111" => color_data <= "000000000000";
      when "010111100001000" => color_data <= "000000000000";
      when "010111100001001" => color_data <= "000000000000";
      when "010111100001010" => color_data <= "000000000000";
      when "010111100001011" => color_data <= "000000000000";
      when "010111100001100" => color_data <= "000000000000";
      when "010111100001101" => color_data <= "000000000000";
      when "010111100001110" => color_data <= "000000000000";
      when "010111100001111" => color_data <= "000000000000";
      when "010111100010000" => color_data <= "000000000000";
      when "010111100010001" => color_data <= "000000000000";
      when "010111100010010" => color_data <= "000000000000";
      when "010111100010011" => color_data <= "000000000000";
      when "010111100010100" => color_data <= "000000000000";
      when "010111100010101" => color_data <= "000000000000";
      when "010111100010110" => color_data <= "000000000000";
      when "010111100010111" => color_data <= "000000000000";
      when "010111100011000" => color_data <= "000000000000";
      when "010111100011001" => color_data <= "000000000000";
      when "010111100011010" => color_data <= "000000000000";
      when "010111100011011" => color_data <= "000000000000";
      when "010111100011100" => color_data <= "000000000000";
      when "010111100011101" => color_data <= "000000000000";
      when "010111100011110" => color_data <= "000000000000";
      when "010111100011111" => color_data <= "000000000000";
      when "010111100100000" => color_data <= "000000000000";
      when "010111100100001" => color_data <= "000000000000";
      when "010111100100010" => color_data <= "000000000000";
      when "010111100100011" => color_data <= "000000000000";
      when "010111100100100" => color_data <= "000000000000";
      when "010111100100101" => color_data <= "000000000000";
      when "010111100100110" => color_data <= "000000000000";
      when "010111100100111" => color_data <= "000000000000";
      when "010111100101000" => color_data <= "000000000000";
      when "010111100101001" => color_data <= "000000000000";
      when "010111100101010" => color_data <= "000000000000";
      when "010111100101011" => color_data <= "000000000000";
      when "010111100101100" => color_data <= "000000000000";
      when "010111100101101" => color_data <= "000000000000";
      when "010111100101110" => color_data <= "001100110010";
      when "010111100101111" => color_data <= "111110110000";
      when "010111100110000" => color_data <= "111111000001";
      when "010111100110001" => color_data <= "111111000001";
      when "010111100110010" => color_data <= "111111000001";
      when "010111100110011" => color_data <= "111111000001";
      when "010111100110100" => color_data <= "111111000001";
      when "010111100110101" => color_data <= "111110110000";
      when "010111100110110" => color_data <= "100001110010";
      when "010111100110111" => color_data <= "000000000000";
      when "010111100111000" => color_data <= "000000000000";
      when "010111100111001" => color_data <= "000000000000";
      when "010111100111010" => color_data <= "000000000000";
      when "010111100111011" => color_data <= "000000000000";
      when "010111100111100" => color_data <= "000000000000";
      when "010111100111101" => color_data <= "000000000000";
      when "010111100111110" => color_data <= "000000000000";
      when "010111100111111" => color_data <= "000000000000";
      when "010111101000000" => color_data <= "000000000000";
      when "010111101000001" => color_data <= "000000000000";
      when "010111101000010" => color_data <= "000000000000";
      when "010111101000011" => color_data <= "000000000000";
      when "010111101000100" => color_data <= "000000000000";
      when "010111101000101" => color_data <= "000000000000";
      when "010111101000110" => color_data <= "000000000000";
      when "010111101000111" => color_data <= "000000000000";
      when "010111101001000" => color_data <= "000000000000";
      when "010111101001001" => color_data <= "000000000000";
      when "010111101001010" => color_data <= "000000000000";
      when "010111101001011" => color_data <= "000000000000";
      when "010111101001100" => color_data <= "000000000000";
      when "010111101001101" => color_data <= "000000000000";
      when "010111101001110" => color_data <= "000000000000";
      when "010111101001111" => color_data <= "000000000000";
      when "010111101010000" => color_data <= "000000000000";
      when "010111101010001" => color_data <= "000000000000";
      when "010111101010010" => color_data <= "000000000000";
      when "010111101010011" => color_data <= "000000000000";
      when "010111101010100" => color_data <= "000000000000";
      when "010111101010101" => color_data <= "000000000000";
      when "010111101010110" => color_data <= "000000000000";
      when "010111101010111" => color_data <= "000000000000";
      when "010111101011000" => color_data <= "000000000000";
      when "010111101011001" => color_data <= "000000000000";
      when "010111101011010" => color_data <= "000000000000";
      when "010111101011011" => color_data <= "000000000000";
      when "010111101011100" => color_data <= "000000000000";
      when "010111101011101" => color_data <= "000000000000";
      when "010111101011110" => color_data <= "000000000000";
      when "010111101011111" => color_data <= "000000000000";
      when "010111101100000" => color_data <= "000000000000";
      when "010111101100001" => color_data <= "000000000000";
      when "010111101100010" => color_data <= "000000000000";
      when "010111101100011" => color_data <= "000000000000";
      when "010111110000000" => color_data <= "000000000000";
      when "010111110000001" => color_data <= "000000000000";
      when "010111110000010" => color_data <= "000000000000";
      when "010111110000011" => color_data <= "000000000000";
      when "010111110000100" => color_data <= "000000000000";
      when "010111110000101" => color_data <= "000000000000";
      when "010111110000110" => color_data <= "000000000000";
      when "010111110000111" => color_data <= "000000000000";
      when "010111110001000" => color_data <= "000000000000";
      when "010111110001001" => color_data <= "000000000000";
      when "010111110001010" => color_data <= "000000000000";
      when "010111110001011" => color_data <= "000000000000";
      when "010111110001100" => color_data <= "000000000000";
      when "010111110001101" => color_data <= "000000000000";
      when "010111110001110" => color_data <= "000000000000";
      when "010111110001111" => color_data <= "000000000000";
      when "010111110010000" => color_data <= "000000000000";
      when "010111110010001" => color_data <= "000000000000";
      when "010111110010010" => color_data <= "000000000000";
      when "010111110010011" => color_data <= "000000000000";
      when "010111110010100" => color_data <= "000000000000";
      when "010111110010101" => color_data <= "000000000000";
      when "010111110010110" => color_data <= "000000000000";
      when "010111110010111" => color_data <= "000000000000";
      when "010111110011000" => color_data <= "000000000000";
      when "010111110011001" => color_data <= "000000000000";
      when "010111110011010" => color_data <= "000000000000";
      when "010111110011011" => color_data <= "000000000000";
      when "010111110011100" => color_data <= "000000000000";
      when "010111110011101" => color_data <= "000000000000";
      when "010111110011110" => color_data <= "000000000000";
      when "010111110011111" => color_data <= "000000000000";
      when "010111110100000" => color_data <= "000000000000";
      when "010111110100001" => color_data <= "000000000000";
      when "010111110100010" => color_data <= "000000000000";
      when "010111110100011" => color_data <= "000000000000";
      when "010111110100100" => color_data <= "000000000000";
      when "010111110100101" => color_data <= "000000000000";
      when "010111110100110" => color_data <= "000000000000";
      when "010111110100111" => color_data <= "000000000000";
      when "010111110101000" => color_data <= "000000000000";
      when "010111110101001" => color_data <= "000000000000";
      when "010111110101010" => color_data <= "000000000000";
      when "010111110101011" => color_data <= "000000000000";
      when "010111110101100" => color_data <= "000000000000";
      when "010111110101101" => color_data <= "000000000000";
      when "010111110101110" => color_data <= "001100110010";
      when "010111110101111" => color_data <= "111110110000";
      when "010111110110000" => color_data <= "111111000001";
      when "010111110110001" => color_data <= "111111000001";
      when "010111110110010" => color_data <= "111111000001";
      when "010111110110011" => color_data <= "111111000001";
      when "010111110110100" => color_data <= "111111000001";
      when "010111110110101" => color_data <= "111110110000";
      when "010111110110110" => color_data <= "100001110010";
      when "010111110110111" => color_data <= "000000000000";
      when "010111110111000" => color_data <= "000000000000";
      when "010111110111001" => color_data <= "000000000000";
      when "010111110111010" => color_data <= "000000000000";
      when "010111110111011" => color_data <= "000000000000";
      when "010111110111100" => color_data <= "000000000000";
      when "010111110111101" => color_data <= "000000000000";
      when "010111110111110" => color_data <= "000000000000";
      when "010111110111111" => color_data <= "000000000000";
      when "010111111000000" => color_data <= "000000000000";
      when "010111111000001" => color_data <= "000000000000";
      when "010111111000010" => color_data <= "000000000000";
      when "010111111000011" => color_data <= "000000000000";
      when "010111111000100" => color_data <= "000000000000";
      when "010111111000101" => color_data <= "000000000000";
      when "010111111000110" => color_data <= "000000000000";
      when "010111111000111" => color_data <= "000000000000";
      when "010111111001000" => color_data <= "000000000000";
      when "010111111001001" => color_data <= "000000000000";
      when "010111111001010" => color_data <= "000000000000";
      when "010111111001011" => color_data <= "000000000000";
      when "010111111001100" => color_data <= "000000000000";
      when "010111111001101" => color_data <= "000000000000";
      when "010111111001110" => color_data <= "000000000000";
      when "010111111001111" => color_data <= "000000000000";
      when "010111111010000" => color_data <= "000000000000";
      when "010111111010001" => color_data <= "000000000000";
      when "010111111010010" => color_data <= "000000000000";
      when "010111111010011" => color_data <= "000000000000";
      when "010111111010100" => color_data <= "000000000000";
      when "010111111010101" => color_data <= "000000000000";
      when "010111111010110" => color_data <= "000000000000";
      when "010111111010111" => color_data <= "000000000000";
      when "010111111011000" => color_data <= "000000000000";
      when "010111111011001" => color_data <= "000000000000";
      when "010111111011010" => color_data <= "000000000000";
      when "010111111011011" => color_data <= "000000000000";
      when "010111111011100" => color_data <= "000000000000";
      when "010111111011101" => color_data <= "000000000000";
      when "010111111011110" => color_data <= "000000000000";
      when "010111111011111" => color_data <= "000000000000";
      when "010111111100000" => color_data <= "000000000000";
      when "010111111100001" => color_data <= "000000000000";
      when "010111111100010" => color_data <= "000000000000";
      when "010111111100011" => color_data <= "000000000000";
      when "011000000000000" => color_data <= "000000000000";
      when "011000000000001" => color_data <= "000000000000";
      when "011000000000010" => color_data <= "000000000000";
      when "011000000000011" => color_data <= "000000000000";
      when "011000000000100" => color_data <= "000000000000";
      when "011000000000101" => color_data <= "000000000000";
      when "011000000000110" => color_data <= "000000000000";
      when "011000000000111" => color_data <= "000000000000";
      when "011000000001000" => color_data <= "000000000000";
      when "011000000001001" => color_data <= "000000000000";
      when "011000000001010" => color_data <= "000000000000";
      when "011000000001011" => color_data <= "000000000000";
      when "011000000001100" => color_data <= "000000000000";
      when "011000000001101" => color_data <= "000000000000";
      when "011000000001110" => color_data <= "000000000000";
      when "011000000001111" => color_data <= "000000000000";
      when "011000000010000" => color_data <= "000000000000";
      when "011000000010001" => color_data <= "000000000000";
      when "011000000010010" => color_data <= "000000000000";
      when "011000000010011" => color_data <= "000000000000";
      when "011000000010100" => color_data <= "000000000000";
      when "011000000010101" => color_data <= "000000000000";
      when "011000000010110" => color_data <= "000000000000";
      when "011000000010111" => color_data <= "000000000000";
      when "011000000011000" => color_data <= "000000000000";
      when "011000000011001" => color_data <= "000000000000";
      when "011000000011010" => color_data <= "000000000000";
      when "011000000011011" => color_data <= "000000000000";
      when "011000000011100" => color_data <= "000000000000";
      when "011000000011101" => color_data <= "000000000000";
      when "011000000011110" => color_data <= "000000000000";
      when "011000000011111" => color_data <= "000000000000";
      when "011000000100000" => color_data <= "000000000000";
      when "011000000100001" => color_data <= "000000000000";
      when "011000000100010" => color_data <= "000000000000";
      when "011000000100011" => color_data <= "000000000000";
      when "011000000100100" => color_data <= "000000000000";
      when "011000000100101" => color_data <= "000000000000";
      when "011000000100110" => color_data <= "000000000000";
      when "011000000100111" => color_data <= "000000000000";
      when "011000000101000" => color_data <= "000000000000";
      when "011000000101001" => color_data <= "000000000000";
      when "011000000101010" => color_data <= "000000000000";
      when "011000000101011" => color_data <= "000000000000";
      when "011000000101100" => color_data <= "000000000000";
      when "011000000101101" => color_data <= "000000000000";
      when "011000000101110" => color_data <= "001100110010";
      when "011000000101111" => color_data <= "111110110000";
      when "011000000110000" => color_data <= "111111000001";
      when "011000000110001" => color_data <= "111111000001";
      when "011000000110010" => color_data <= "111111000001";
      when "011000000110011" => color_data <= "111111000001";
      when "011000000110100" => color_data <= "111111000001";
      when "011000000110101" => color_data <= "111110110000";
      when "011000000110110" => color_data <= "100001110010";
      when "011000000110111" => color_data <= "000000000000";
      when "011000000111000" => color_data <= "000000000000";
      when "011000000111001" => color_data <= "000000000000";
      when "011000000111010" => color_data <= "000000000000";
      when "011000000111011" => color_data <= "000000000000";
      when "011000000111100" => color_data <= "000000000000";
      when "011000000111101" => color_data <= "000000000000";
      when "011000000111110" => color_data <= "000000000000";
      when "011000000111111" => color_data <= "000000000000";
      when "011000001000000" => color_data <= "000000000000";
      when "011000001000001" => color_data <= "000000000000";
      when "011000001000010" => color_data <= "000000000000";
      when "011000001000011" => color_data <= "000000000000";
      when "011000001000100" => color_data <= "000000000000";
      when "011000001000101" => color_data <= "000000000000";
      when "011000001000110" => color_data <= "000000000000";
      when "011000001000111" => color_data <= "000000000000";
      when "011000001001000" => color_data <= "000000000000";
      when "011000001001001" => color_data <= "000000000000";
      when "011000001001010" => color_data <= "000000000000";
      when "011000001001011" => color_data <= "000000000000";
      when "011000001001100" => color_data <= "000000000000";
      when "011000001001101" => color_data <= "000000000000";
      when "011000001001110" => color_data <= "000000000000";
      when "011000001001111" => color_data <= "000000000000";
      when "011000001010000" => color_data <= "000000000000";
      when "011000001010001" => color_data <= "000000000000";
      when "011000001010010" => color_data <= "000000000000";
      when "011000001010011" => color_data <= "000000000000";
      when "011000001010100" => color_data <= "000000000000";
      when "011000001010101" => color_data <= "000000000000";
      when "011000001010110" => color_data <= "000000000000";
      when "011000001010111" => color_data <= "000000000000";
      when "011000001011000" => color_data <= "000000000000";
      when "011000001011001" => color_data <= "000000000000";
      when "011000001011010" => color_data <= "000000000000";
      when "011000001011011" => color_data <= "000000000000";
      when "011000001011100" => color_data <= "000000000000";
      when "011000001011101" => color_data <= "000000000000";
      when "011000001011110" => color_data <= "000000000000";
      when "011000001011111" => color_data <= "000000000000";
      when "011000001100000" => color_data <= "000000000000";
      when "011000001100001" => color_data <= "000000000000";
      when "011000001100010" => color_data <= "000000000000";
      when "011000001100011" => color_data <= "000000000000";
      when "011000010000000" => color_data <= "000000000000";
      when "011000010000001" => color_data <= "000000000000";
      when "011000010000010" => color_data <= "000000000000";
      when "011000010000011" => color_data <= "000000000000";
      when "011000010000100" => color_data <= "000000000000";
      when "011000010000101" => color_data <= "000000000000";
      when "011000010000110" => color_data <= "000000000000";
      when "011000010000111" => color_data <= "000000000000";
      when "011000010001000" => color_data <= "000000000000";
      when "011000010001001" => color_data <= "000000000000";
      when "011000010001010" => color_data <= "000000000000";
      when "011000010001011" => color_data <= "000000000000";
      when "011000010001100" => color_data <= "000000000000";
      when "011000010001101" => color_data <= "000000000000";
      when "011000010001110" => color_data <= "000000000000";
      when "011000010001111" => color_data <= "000000000000";
      when "011000010010000" => color_data <= "000000000000";
      when "011000010010001" => color_data <= "000000000000";
      when "011000010010010" => color_data <= "000000000000";
      when "011000010010011" => color_data <= "000000000000";
      when "011000010010100" => color_data <= "000000000000";
      when "011000010010101" => color_data <= "000000000000";
      when "011000010010110" => color_data <= "000000000000";
      when "011000010010111" => color_data <= "000000000000";
      when "011000010011000" => color_data <= "000000000000";
      when "011000010011001" => color_data <= "000000000000";
      when "011000010011010" => color_data <= "000000000000";
      when "011000010011011" => color_data <= "000000000000";
      when "011000010011100" => color_data <= "000000000000";
      when "011000010011101" => color_data <= "000000000000";
      when "011000010011110" => color_data <= "000000000000";
      when "011000010011111" => color_data <= "000000000000";
      when "011000010100000" => color_data <= "000000000000";
      when "011000010100001" => color_data <= "000000000000";
      when "011000010100010" => color_data <= "000000000000";
      when "011000010100011" => color_data <= "000000000000";
      when "011000010100100" => color_data <= "000000000000";
      when "011000010100101" => color_data <= "000000000000";
      when "011000010100110" => color_data <= "000000000000";
      when "011000010100111" => color_data <= "000000000000";
      when "011000010101000" => color_data <= "000000000000";
      when "011000010101001" => color_data <= "000000000000";
      when "011000010101010" => color_data <= "000000000000";
      when "011000010101011" => color_data <= "000000000000";
      when "011000010101100" => color_data <= "000000000000";
      when "011000010101101" => color_data <= "000000000000";
      when "011000010101110" => color_data <= "001100110010";
      when "011000010101111" => color_data <= "111110110000";
      when "011000010110000" => color_data <= "111111000001";
      when "011000010110001" => color_data <= "111111000001";
      when "011000010110010" => color_data <= "111111000001";
      when "011000010110011" => color_data <= "111111000001";
      when "011000010110100" => color_data <= "111111000001";
      when "011000010110101" => color_data <= "111110110000";
      when "011000010110110" => color_data <= "100001110010";
      when "011000010110111" => color_data <= "000000000000";
      when "011000010111000" => color_data <= "000000000000";
      when "011000010111001" => color_data <= "000000000000";
      when "011000010111010" => color_data <= "000000000000";
      when "011000010111011" => color_data <= "000000000000";
      when "011000010111100" => color_data <= "000000000000";
      when "011000010111101" => color_data <= "000000000000";
      when "011000010111110" => color_data <= "000000000000";
      when "011000010111111" => color_data <= "000000000000";
      when "011000011000000" => color_data <= "000000000000";
      when "011000011000001" => color_data <= "000000000000";
      when "011000011000010" => color_data <= "000000000000";
      when "011000011000011" => color_data <= "000000000000";
      when "011000011000100" => color_data <= "000000000000";
      when "011000011000101" => color_data <= "000000000000";
      when "011000011000110" => color_data <= "000000000000";
      when "011000011000111" => color_data <= "000000000000";
      when "011000011001000" => color_data <= "000000000000";
      when "011000011001001" => color_data <= "000000000000";
      when "011000011001010" => color_data <= "000000000000";
      when "011000011001011" => color_data <= "000000000000";
      when "011000011001100" => color_data <= "000000000000";
      when "011000011001101" => color_data <= "000000000000";
      when "011000011001110" => color_data <= "000000000000";
      when "011000011001111" => color_data <= "000000000000";
      when "011000011010000" => color_data <= "000000000000";
      when "011000011010001" => color_data <= "000000000000";
      when "011000011010010" => color_data <= "000000000000";
      when "011000011010011" => color_data <= "000000000000";
      when "011000011010100" => color_data <= "000000000000";
      when "011000011010101" => color_data <= "000000000000";
      when "011000011010110" => color_data <= "000000000000";
      when "011000011010111" => color_data <= "000000000000";
      when "011000011011000" => color_data <= "000000000000";
      when "011000011011001" => color_data <= "000000000000";
      when "011000011011010" => color_data <= "000000000000";
      when "011000011011011" => color_data <= "000000000000";
      when "011000011011100" => color_data <= "000000000000";
      when "011000011011101" => color_data <= "000000000000";
      when "011000011011110" => color_data <= "000000000000";
      when "011000011011111" => color_data <= "000000000000";
      when "011000011100000" => color_data <= "000000000000";
      when "011000011100001" => color_data <= "000000000000";
      when "011000011100010" => color_data <= "000000000000";
      when "011000011100011" => color_data <= "000000000000";
      when "011000100000000" => color_data <= "000000000000";
      when "011000100000001" => color_data <= "000000000000";
      when "011000100000010" => color_data <= "000000000000";
      when "011000100000011" => color_data <= "000000000000";
      when "011000100000100" => color_data <= "000000000000";
      when "011000100000101" => color_data <= "000000000000";
      when "011000100000110" => color_data <= "000000000000";
      when "011000100000111" => color_data <= "000000000000";
      when "011000100001000" => color_data <= "000000000000";
      when "011000100001001" => color_data <= "000000000000";
      when "011000100001010" => color_data <= "000000000000";
      when "011000100001011" => color_data <= "000000000000";
      when "011000100001100" => color_data <= "000000000000";
      when "011000100001101" => color_data <= "000000000000";
      when "011000100001110" => color_data <= "000000000000";
      when "011000100001111" => color_data <= "000000000000";
      when "011000100010000" => color_data <= "000000000000";
      when "011000100010001" => color_data <= "000000000000";
      when "011000100010010" => color_data <= "000000000000";
      when "011000100010011" => color_data <= "000000000000";
      when "011000100010100" => color_data <= "000000000000";
      when "011000100010101" => color_data <= "000000000000";
      when "011000100010110" => color_data <= "000000000000";
      when "011000100010111" => color_data <= "000000000000";
      when "011000100011000" => color_data <= "000000000000";
      when "011000100011001" => color_data <= "000000000000";
      when "011000100011010" => color_data <= "000000000000";
      when "011000100011011" => color_data <= "000000000000";
      when "011000100011100" => color_data <= "000000000000";
      when "011000100011101" => color_data <= "000000000000";
      when "011000100011110" => color_data <= "000000000000";
      when "011000100011111" => color_data <= "000000000000";
      when "011000100100000" => color_data <= "000000000000";
      when "011000100100001" => color_data <= "000000000000";
      when "011000100100010" => color_data <= "000000000000";
      when "011000100100011" => color_data <= "000000000000";
      when "011000100100100" => color_data <= "000000000000";
      when "011000100100101" => color_data <= "000000000000";
      when "011000100100110" => color_data <= "000000000000";
      when "011000100100111" => color_data <= "000000000000";
      when "011000100101000" => color_data <= "000000000000";
      when "011000100101001" => color_data <= "000000000000";
      when "011000100101010" => color_data <= "000000000000";
      when "011000100101011" => color_data <= "000000000000";
      when "011000100101100" => color_data <= "000000000000";
      when "011000100101101" => color_data <= "000000000000";
      when "011000100101110" => color_data <= "001100110010";
      when "011000100101111" => color_data <= "111110110000";
      when "011000100110000" => color_data <= "111111000001";
      when "011000100110001" => color_data <= "111111000001";
      when "011000100110010" => color_data <= "111111000001";
      when "011000100110011" => color_data <= "111111000001";
      when "011000100110100" => color_data <= "111111000001";
      when "011000100110101" => color_data <= "111110110000";
      when "011000100110110" => color_data <= "100001110010";
      when "011000100110111" => color_data <= "000000000000";
      when "011000100111000" => color_data <= "000000000000";
      when "011000100111001" => color_data <= "000000000000";
      when "011000100111010" => color_data <= "000000000000";
      when "011000100111011" => color_data <= "000000000000";
      when "011000100111100" => color_data <= "000000000000";
      when "011000100111101" => color_data <= "000000000000";
      when "011000100111110" => color_data <= "000000000000";
      when "011000100111111" => color_data <= "000000000000";
      when "011000101000000" => color_data <= "000000000000";
      when "011000101000001" => color_data <= "000000000000";
      when "011000101000010" => color_data <= "000000000000";
      when "011000101000011" => color_data <= "000000000000";
      when "011000101000100" => color_data <= "000000000000";
      when "011000101000101" => color_data <= "000000000000";
      when "011000101000110" => color_data <= "000000000000";
      when "011000101000111" => color_data <= "000000000000";
      when "011000101001000" => color_data <= "000000000000";
      when "011000101001001" => color_data <= "000000000000";
      when "011000101001010" => color_data <= "000000000000";
      when "011000101001011" => color_data <= "000000000000";
      when "011000101001100" => color_data <= "000000000000";
      when "011000101001101" => color_data <= "000000000000";
      when "011000101001110" => color_data <= "000000000000";
      when "011000101001111" => color_data <= "000000000000";
      when "011000101010000" => color_data <= "000000000000";
      when "011000101010001" => color_data <= "000000000000";
      when "011000101010010" => color_data <= "000000000000";
      when "011000101010011" => color_data <= "000000000000";
      when "011000101010100" => color_data <= "000000000000";
      when "011000101010101" => color_data <= "000000000000";
      when "011000101010110" => color_data <= "000000000000";
      when "011000101010111" => color_data <= "000000000000";
      when "011000101011000" => color_data <= "000000000000";
      when "011000101011001" => color_data <= "000000000000";
      when "011000101011010" => color_data <= "000000000000";
      when "011000101011011" => color_data <= "000000000000";
      when "011000101011100" => color_data <= "000000000000";
      when "011000101011101" => color_data <= "000000000000";
      when "011000101011110" => color_data <= "000000000000";
      when "011000101011111" => color_data <= "000000000000";
      when "011000101100000" => color_data <= "000000000000";
      when "011000101100001" => color_data <= "000000000000";
      when "011000101100010" => color_data <= "000000000000";
      when "011000101100011" => color_data <= "000000000000";
      when "011000110000000" => color_data <= "000000000000";
      when "011000110000001" => color_data <= "000000000000";
      when "011000110000010" => color_data <= "000000000000";
      when "011000110000011" => color_data <= "000000000000";
      when "011000110000100" => color_data <= "000000000000";
      when "011000110000101" => color_data <= "000000000000";
      when "011000110000110" => color_data <= "000000000000";
      when "011000110000111" => color_data <= "000000000000";
      when "011000110001000" => color_data <= "000000000000";
      when "011000110001001" => color_data <= "000000000000";
      when "011000110001010" => color_data <= "000000000000";
      when "011000110001011" => color_data <= "000000000000";
      when "011000110001100" => color_data <= "000000000000";
      when "011000110001101" => color_data <= "000000000000";
      when "011000110001110" => color_data <= "000000000000";
      when "011000110001111" => color_data <= "000000000000";
      when "011000110010000" => color_data <= "000000000000";
      when "011000110010001" => color_data <= "000000000000";
      when "011000110010010" => color_data <= "000000000000";
      when "011000110010011" => color_data <= "000000000000";
      when "011000110010100" => color_data <= "000000000000";
      when "011000110010101" => color_data <= "000000000000";
      when "011000110010110" => color_data <= "000000000000";
      when "011000110010111" => color_data <= "000000000000";
      when "011000110011000" => color_data <= "000000000000";
      when "011000110011001" => color_data <= "000000000000";
      when "011000110011010" => color_data <= "000000000000";
      when "011000110011011" => color_data <= "000000000000";
      when "011000110011100" => color_data <= "000000000000";
      when "011000110011101" => color_data <= "000000000000";
      when "011000110011110" => color_data <= "000000000000";
      when "011000110011111" => color_data <= "000000000000";
      when "011000110100000" => color_data <= "000000000000";
      when "011000110100001" => color_data <= "000000000000";
      when "011000110100010" => color_data <= "000000000000";
      when "011000110100011" => color_data <= "000000000000";
      when "011000110100100" => color_data <= "000000000000";
      when "011000110100101" => color_data <= "000000000000";
      when "011000110100110" => color_data <= "000000000000";
      when "011000110100111" => color_data <= "000000000000";
      when "011000110101000" => color_data <= "000000000000";
      when "011000110101001" => color_data <= "000000000000";
      when "011000110101010" => color_data <= "000000000000";
      when "011000110101011" => color_data <= "000000000000";
      when "011000110101100" => color_data <= "000000000000";
      when "011000110101101" => color_data <= "000000000000";
      when "011000110101110" => color_data <= "010000110010";
      when "011000110101111" => color_data <= "111110110000";
      when "011000110110000" => color_data <= "111111000001";
      when "011000110110001" => color_data <= "111111000001";
      when "011000110110010" => color_data <= "111111000001";
      when "011000110110011" => color_data <= "111111000001";
      when "011000110110100" => color_data <= "111111000001";
      when "011000110110101" => color_data <= "111110110000";
      when "011000110110110" => color_data <= "100001110010";
      when "011000110110111" => color_data <= "000000000000";
      when "011000110111000" => color_data <= "000000000000";
      when "011000110111001" => color_data <= "000000000000";
      when "011000110111010" => color_data <= "000000000000";
      when "011000110111011" => color_data <= "000000000000";
      when "011000110111100" => color_data <= "000000000000";
      when "011000110111101" => color_data <= "000000000000";
      when "011000110111110" => color_data <= "000000000000";
      when "011000110111111" => color_data <= "000000000000";
      when "011000111000000" => color_data <= "000000000000";
      when "011000111000001" => color_data <= "000000000000";
      when "011000111000010" => color_data <= "000000000000";
      when "011000111000011" => color_data <= "000000000000";
      when "011000111000100" => color_data <= "000000000000";
      when "011000111000101" => color_data <= "000000000000";
      when "011000111000110" => color_data <= "000000000000";
      when "011000111000111" => color_data <= "000000000000";
      when "011000111001000" => color_data <= "000000000000";
      when "011000111001001" => color_data <= "000000000000";
      when "011000111001010" => color_data <= "000000000000";
      when "011000111001011" => color_data <= "000000000000";
      when "011000111001100" => color_data <= "000000000000";
      when "011000111001101" => color_data <= "000000000000";
      when "011000111001110" => color_data <= "000000000000";
      when "011000111001111" => color_data <= "000000000000";
      when "011000111010000" => color_data <= "000000000000";
      when "011000111010001" => color_data <= "000000000000";
      when "011000111010010" => color_data <= "000000000000";
      when "011000111010011" => color_data <= "000000000000";
      when "011000111010100" => color_data <= "000000000000";
      when "011000111010101" => color_data <= "000000000000";
      when "011000111010110" => color_data <= "000000000000";
      when "011000111010111" => color_data <= "000000000000";
      when "011000111011000" => color_data <= "000000000000";
      when "011000111011001" => color_data <= "000000000000";
      when "011000111011010" => color_data <= "000000000000";
      when "011000111011011" => color_data <= "000000000000";
      when "011000111011100" => color_data <= "000000000000";
      when "011000111011101" => color_data <= "000000000000";
      when "011000111011110" => color_data <= "000000000000";
      when "011000111011111" => color_data <= "000000000000";
      when "011000111100000" => color_data <= "000000000000";
      when "011000111100001" => color_data <= "000000000000";
      when "011000111100010" => color_data <= "000000000000";
      when "011000111100011" => color_data <= "000000000000";
      when "011001000000000" => color_data <= "000000000000";
      when "011001000000001" => color_data <= "000000000000";
      when "011001000000010" => color_data <= "000000000000";
      when "011001000000011" => color_data <= "000000000000";
      when "011001000000100" => color_data <= "000000000000";
      when "011001000000101" => color_data <= "000000000000";
      when "011001000000110" => color_data <= "000000000000";
      when "011001000000111" => color_data <= "000000000000";
      when "011001000001000" => color_data <= "000000000000";
      when "011001000001001" => color_data <= "000000000000";
      when "011001000001010" => color_data <= "000000000000";
      when "011001000001011" => color_data <= "000000000000";
      when "011001000001100" => color_data <= "000000000000";
      when "011001000001101" => color_data <= "000000000000";
      when "011001000001110" => color_data <= "000000000000";
      when "011001000001111" => color_data <= "000000000000";
      when "011001000010000" => color_data <= "000000000000";
      when "011001000010001" => color_data <= "000000000000";
      when "011001000010010" => color_data <= "000000000000";
      when "011001000010011" => color_data <= "000000000000";
      when "011001000010100" => color_data <= "000000000000";
      when "011001000010101" => color_data <= "000000000000";
      when "011001000010110" => color_data <= "000000000000";
      when "011001000010111" => color_data <= "000000000000";
      when "011001000011000" => color_data <= "000000000000";
      when "011001000011001" => color_data <= "000000000000";
      when "011001000011010" => color_data <= "000000000000";
      when "011001000011011" => color_data <= "000000000000";
      when "011001000011100" => color_data <= "000000000000";
      when "011001000011101" => color_data <= "000000000000";
      when "011001000011110" => color_data <= "000000000000";
      when "011001000011111" => color_data <= "000000000000";
      when "011001000100000" => color_data <= "000000000000";
      when "011001000100001" => color_data <= "000000000000";
      when "011001000100010" => color_data <= "000000000000";
      when "011001000100011" => color_data <= "000000000000";
      when "011001000100100" => color_data <= "000000000000";
      when "011001000100101" => color_data <= "000000000000";
      when "011001000100110" => color_data <= "000000000000";
      when "011001000100111" => color_data <= "000000000000";
      when "011001000101000" => color_data <= "000000000000";
      when "011001000101001" => color_data <= "000000000000";
      when "011001000101010" => color_data <= "000000000000";
      when "011001000101011" => color_data <= "000000000000";
      when "011001000101100" => color_data <= "000000000000";
      when "011001000101101" => color_data <= "000000000000";
      when "011001000101110" => color_data <= "010000110010";
      when "011001000101111" => color_data <= "111110110000";
      when "011001000110000" => color_data <= "111111000001";
      when "011001000110001" => color_data <= "111111000001";
      when "011001000110010" => color_data <= "111111000001";
      when "011001000110011" => color_data <= "111111000001";
      when "011001000110100" => color_data <= "111111000001";
      when "011001000110101" => color_data <= "111110110000";
      when "011001000110110" => color_data <= "100001110010";
      when "011001000110111" => color_data <= "000000000000";
      when "011001000111000" => color_data <= "000000000000";
      when "011001000111001" => color_data <= "000000000000";
      when "011001000111010" => color_data <= "000000000000";
      when "011001000111011" => color_data <= "000000000000";
      when "011001000111100" => color_data <= "000000000000";
      when "011001000111101" => color_data <= "000000000000";
      when "011001000111110" => color_data <= "000000000000";
      when "011001000111111" => color_data <= "000000000000";
      when "011001001000000" => color_data <= "000000000000";
      when "011001001000001" => color_data <= "000000000000";
      when "011001001000010" => color_data <= "000000000000";
      when "011001001000011" => color_data <= "000000000000";
      when "011001001000100" => color_data <= "000000000000";
      when "011001001000101" => color_data <= "000000000000";
      when "011001001000110" => color_data <= "000000000000";
      when "011001001000111" => color_data <= "000000000000";
      when "011001001001000" => color_data <= "000000000000";
      when "011001001001001" => color_data <= "000000000000";
      when "011001001001010" => color_data <= "000000000000";
      when "011001001001011" => color_data <= "000000000000";
      when "011001001001100" => color_data <= "000000000000";
      when "011001001001101" => color_data <= "000000000000";
      when "011001001001110" => color_data <= "000000000000";
      when "011001001001111" => color_data <= "000000000000";
      when "011001001010000" => color_data <= "000000000000";
      when "011001001010001" => color_data <= "000000000000";
      when "011001001010010" => color_data <= "000000000000";
      when "011001001010011" => color_data <= "000000000000";
      when "011001001010100" => color_data <= "000000000000";
      when "011001001010101" => color_data <= "000000000000";
      when "011001001010110" => color_data <= "000000000000";
      when "011001001010111" => color_data <= "000000000000";
      when "011001001011000" => color_data <= "000000000000";
      when "011001001011001" => color_data <= "000000000000";
      when "011001001011010" => color_data <= "000000000000";
      when "011001001011011" => color_data <= "000000000000";
      when "011001001011100" => color_data <= "000000000000";
      when "011001001011101" => color_data <= "000000000000";
      when "011001001011110" => color_data <= "000000000000";
      when "011001001011111" => color_data <= "000000000000";
      when "011001001100000" => color_data <= "000000000000";
      when "011001001100001" => color_data <= "000000000000";
      when "011001001100010" => color_data <= "000000000000";
      when "011001001100011" => color_data <= "000000000000";
      when "011001010000000" => color_data <= "000000000000";
      when "011001010000001" => color_data <= "000000000000";
      when "011001010000010" => color_data <= "000000000000";
      when "011001010000011" => color_data <= "000000000000";
      when "011001010000100" => color_data <= "000000000000";
      when "011001010000101" => color_data <= "000000000000";
      when "011001010000110" => color_data <= "000000000000";
      when "011001010000111" => color_data <= "000000000000";
      when "011001010001000" => color_data <= "000000000000";
      when "011001010001001" => color_data <= "000000000000";
      when "011001010001010" => color_data <= "000000000000";
      when "011001010001011" => color_data <= "000000000000";
      when "011001010001100" => color_data <= "000000000000";
      when "011001010001101" => color_data <= "000000000000";
      when "011001010001110" => color_data <= "000000000000";
      when "011001010001111" => color_data <= "000000000000";
      when "011001010010000" => color_data <= "000000000000";
      when "011001010010001" => color_data <= "000000000000";
      when "011001010010010" => color_data <= "000000000000";
      when "011001010010011" => color_data <= "000000000000";
      when "011001010010100" => color_data <= "000000000000";
      when "011001010010101" => color_data <= "000000000000";
      when "011001010010110" => color_data <= "000000000000";
      when "011001010010111" => color_data <= "000000000000";
      when "011001010011000" => color_data <= "000000000000";
      when "011001010011001" => color_data <= "000000000000";
      when "011001010011010" => color_data <= "000000000000";
      when "011001010011011" => color_data <= "000000000000";
      when "011001010011100" => color_data <= "000000000000";
      when "011001010011101" => color_data <= "000000000000";
      when "011001010011110" => color_data <= "000000000000";
      when "011001010011111" => color_data <= "000000000000";
      when "011001010100000" => color_data <= "000000000000";
      when "011001010100001" => color_data <= "000000000000";
      when "011001010100010" => color_data <= "000000000000";
      when "011001010100011" => color_data <= "000000000000";
      when "011001010100100" => color_data <= "000000000000";
      when "011001010100101" => color_data <= "000000000000";
      when "011001010100110" => color_data <= "000000000000";
      when "011001010100111" => color_data <= "000000000000";
      when "011001010101000" => color_data <= "000000000000";
      when "011001010101001" => color_data <= "000000000000";
      when "011001010101010" => color_data <= "000000000000";
      when "011001010101011" => color_data <= "000000000000";
      when "011001010101100" => color_data <= "000000000000";
      when "011001010101101" => color_data <= "000000000000";
      when "011001010101110" => color_data <= "010001000010";
      when "011001010101111" => color_data <= "111110110000";
      when "011001010110000" => color_data <= "111111000001";
      when "011001010110001" => color_data <= "111111000001";
      when "011001010110010" => color_data <= "111111000001";
      when "011001010110011" => color_data <= "111111000001";
      when "011001010110100" => color_data <= "111111000001";
      when "011001010110101" => color_data <= "111110110000";
      when "011001010110110" => color_data <= "100101110010";
      when "011001010110111" => color_data <= "000000000000";
      when "011001010111000" => color_data <= "000000000000";
      when "011001010111001" => color_data <= "000000000000";
      when "011001010111010" => color_data <= "000000000000";
      when "011001010111011" => color_data <= "000000000000";
      when "011001010111100" => color_data <= "000000000000";
      when "011001010111101" => color_data <= "000000000000";
      when "011001010111110" => color_data <= "000000000000";
      when "011001010111111" => color_data <= "000000000000";
      when "011001011000000" => color_data <= "000000000000";
      when "011001011000001" => color_data <= "000000000000";
      when "011001011000010" => color_data <= "000000000000";
      when "011001011000011" => color_data <= "000000000000";
      when "011001011000100" => color_data <= "000000000000";
      when "011001011000101" => color_data <= "000000000000";
      when "011001011000110" => color_data <= "000000000000";
      when "011001011000111" => color_data <= "000000000000";
      when "011001011001000" => color_data <= "000000000000";
      when "011001011001001" => color_data <= "000000000000";
      when "011001011001010" => color_data <= "000000000000";
      when "011001011001011" => color_data <= "000000000000";
      when "011001011001100" => color_data <= "000000000000";
      when "011001011001101" => color_data <= "000000000000";
      when "011001011001110" => color_data <= "000000000000";
      when "011001011001111" => color_data <= "000000000000";
      when "011001011010000" => color_data <= "000000000000";
      when "011001011010001" => color_data <= "000000000000";
      when "011001011010010" => color_data <= "000000000000";
      when "011001011010011" => color_data <= "000000000000";
      when "011001011010100" => color_data <= "000000000000";
      when "011001011010101" => color_data <= "000000000000";
      when "011001011010110" => color_data <= "000000000000";
      when "011001011010111" => color_data <= "000000000000";
      when "011001011011000" => color_data <= "000000000000";
      when "011001011011001" => color_data <= "000000000000";
      when "011001011011010" => color_data <= "000000000000";
      when "011001011011011" => color_data <= "000000000000";
      when "011001011011100" => color_data <= "000000000000";
      when "011001011011101" => color_data <= "000000000000";
      when "011001011011110" => color_data <= "000000000000";
      when "011001011011111" => color_data <= "000000000000";
      when "011001011100000" => color_data <= "000000000000";
      when "011001011100001" => color_data <= "000000000000";
      when "011001011100010" => color_data <= "000000000000";
      when "011001011100011" => color_data <= "000000000000";
      when "011001100000000" => color_data <= "000000000000";
      when "011001100000001" => color_data <= "000000000000";
      when "011001100000010" => color_data <= "000000000000";
      when "011001100000011" => color_data <= "000000000000";
      when "011001100000100" => color_data <= "000000000000";
      when "011001100000101" => color_data <= "000000000000";
      when "011001100000110" => color_data <= "000000000000";
      when "011001100000111" => color_data <= "000000000000";
      when "011001100001000" => color_data <= "000000000000";
      when "011001100001001" => color_data <= "000000000000";
      when "011001100001010" => color_data <= "000000000000";
      when "011001100001011" => color_data <= "000000000000";
      when "011001100001100" => color_data <= "000000000000";
      when "011001100001101" => color_data <= "000000000000";
      when "011001100001110" => color_data <= "000000000000";
      when "011001100001111" => color_data <= "000000000000";
      when "011001100010000" => color_data <= "000000000000";
      when "011001100010001" => color_data <= "000000000000";
      when "011001100010010" => color_data <= "000000000000";
      when "011001100010011" => color_data <= "000000000000";
      when "011001100010100" => color_data <= "000000000000";
      when "011001100010101" => color_data <= "000000000000";
      when "011001100010110" => color_data <= "000000000000";
      when "011001100010111" => color_data <= "000000000000";
      when "011001100011000" => color_data <= "000000000000";
      when "011001100011001" => color_data <= "000000000000";
      when "011001100011010" => color_data <= "000000000000";
      when "011001100011011" => color_data <= "000000000000";
      when "011001100011100" => color_data <= "000000000000";
      when "011001100011101" => color_data <= "000000000000";
      when "011001100011110" => color_data <= "000000000000";
      when "011001100011111" => color_data <= "000000000000";
      when "011001100100000" => color_data <= "000000000000";
      when "011001100100001" => color_data <= "000000000000";
      when "011001100100010" => color_data <= "000000000000";
      when "011001100100011" => color_data <= "000000000000";
      when "011001100100100" => color_data <= "000000000000";
      when "011001100100101" => color_data <= "000000000000";
      when "011001100100110" => color_data <= "000000000000";
      when "011001100100111" => color_data <= "000000000000";
      when "011001100101000" => color_data <= "000000000000";
      when "011001100101001" => color_data <= "000000000000";
      when "011001100101010" => color_data <= "000000000000";
      when "011001100101011" => color_data <= "000000000000";
      when "011001100101100" => color_data <= "000000000000";
      when "011001100101101" => color_data <= "000000000000";
      when "011001100101110" => color_data <= "010101000010";
      when "011001100101111" => color_data <= "111110110000";
      when "011001100110000" => color_data <= "111111000001";
      when "011001100110001" => color_data <= "111111000001";
      when "011001100110010" => color_data <= "111111000001";
      when "011001100110011" => color_data <= "111111000001";
      when "011001100110100" => color_data <= "111111000001";
      when "011001100110101" => color_data <= "111110110000";
      when "011001100110110" => color_data <= "100110000010";
      when "011001100110111" => color_data <= "000000000000";
      when "011001100111000" => color_data <= "000000000000";
      when "011001100111001" => color_data <= "000000000000";
      when "011001100111010" => color_data <= "000000000000";
      when "011001100111011" => color_data <= "000000000000";
      when "011001100111100" => color_data <= "000000000000";
      when "011001100111101" => color_data <= "000000000000";
      when "011001100111110" => color_data <= "000000000000";
      when "011001100111111" => color_data <= "000000000000";
      when "011001101000000" => color_data <= "000000000000";
      when "011001101000001" => color_data <= "000000000000";
      when "011001101000010" => color_data <= "000000000000";
      when "011001101000011" => color_data <= "000000000000";
      when "011001101000100" => color_data <= "000000000000";
      when "011001101000101" => color_data <= "000000000000";
      when "011001101000110" => color_data <= "000000000000";
      when "011001101000111" => color_data <= "000000000000";
      when "011001101001000" => color_data <= "000000000000";
      when "011001101001001" => color_data <= "000000000000";
      when "011001101001010" => color_data <= "000000000000";
      when "011001101001011" => color_data <= "000000000000";
      when "011001101001100" => color_data <= "000000000000";
      when "011001101001101" => color_data <= "000000000000";
      when "011001101001110" => color_data <= "000000000000";
      when "011001101001111" => color_data <= "000000000000";
      when "011001101010000" => color_data <= "000000000000";
      when "011001101010001" => color_data <= "000000000000";
      when "011001101010010" => color_data <= "000000000000";
      when "011001101010011" => color_data <= "000000000000";
      when "011001101010100" => color_data <= "000000000000";
      when "011001101010101" => color_data <= "000000000000";
      when "011001101010110" => color_data <= "000000000000";
      when "011001101010111" => color_data <= "000000000000";
      when "011001101011000" => color_data <= "000000000000";
      when "011001101011001" => color_data <= "000000000000";
      when "011001101011010" => color_data <= "000000000000";
      when "011001101011011" => color_data <= "000000000000";
      when "011001101011100" => color_data <= "000000000000";
      when "011001101011101" => color_data <= "000000000000";
      when "011001101011110" => color_data <= "000000000000";
      when "011001101011111" => color_data <= "000000000000";
      when "011001101100000" => color_data <= "000000000000";
      when "011001101100001" => color_data <= "000000000000";
      when "011001101100010" => color_data <= "000000000000";
      when "011001101100011" => color_data <= "000000000000";
      when "011001110000000" => color_data <= "000000000000";
      when "011001110000001" => color_data <= "000000000000";
      when "011001110000010" => color_data <= "000000000000";
      when "011001110000011" => color_data <= "000000000000";
      when "011001110000100" => color_data <= "000000000000";
      when "011001110000101" => color_data <= "000000000000";
      when "011001110000110" => color_data <= "000000000000";
      when "011001110000111" => color_data <= "000000000000";
      when "011001110001000" => color_data <= "000000000000";
      when "011001110001001" => color_data <= "000000000000";
      when "011001110001010" => color_data <= "000000000000";
      when "011001110001011" => color_data <= "000000000000";
      when "011001110001100" => color_data <= "000000000000";
      when "011001110001101" => color_data <= "000000000000";
      when "011001110001110" => color_data <= "000000000000";
      when "011001110001111" => color_data <= "000000000000";
      when "011001110010000" => color_data <= "000000000000";
      when "011001110010001" => color_data <= "000000000000";
      when "011001110010010" => color_data <= "000000000000";
      when "011001110010011" => color_data <= "000000000000";
      when "011001110010100" => color_data <= "000000000000";
      when "011001110010101" => color_data <= "000000000000";
      when "011001110010110" => color_data <= "000000000000";
      when "011001110010111" => color_data <= "000000000000";
      when "011001110011000" => color_data <= "000000000000";
      when "011001110011001" => color_data <= "000000000000";
      when "011001110011010" => color_data <= "000000000000";
      when "011001110011011" => color_data <= "000000000000";
      when "011001110011100" => color_data <= "000000000000";
      when "011001110011101" => color_data <= "000000000000";
      when "011001110011110" => color_data <= "000000000000";
      when "011001110011111" => color_data <= "000000000000";
      when "011001110100000" => color_data <= "000000000000";
      when "011001110100001" => color_data <= "000000000000";
      when "011001110100010" => color_data <= "000000000000";
      when "011001110100011" => color_data <= "000000000000";
      when "011001110100100" => color_data <= "000000000000";
      when "011001110100101" => color_data <= "000000000000";
      when "011001110100110" => color_data <= "000000000000";
      when "011001110100111" => color_data <= "000000000000";
      when "011001110101000" => color_data <= "000000000000";
      when "011001110101001" => color_data <= "000000000000";
      when "011001110101010" => color_data <= "000000000000";
      when "011001110101011" => color_data <= "000000000000";
      when "011001110101100" => color_data <= "000000000000";
      when "011001110101101" => color_data <= "000000000000";
      when "011001110101110" => color_data <= "011001010011";
      when "011001110101111" => color_data <= "111110110000";
      when "011001110110000" => color_data <= "111111000001";
      when "011001110110001" => color_data <= "111111000001";
      when "011001110110010" => color_data <= "111111000001";
      when "011001110110011" => color_data <= "111111000001";
      when "011001110110100" => color_data <= "111111000001";
      when "011001110110101" => color_data <= "111110110000";
      when "011001110110110" => color_data <= "101010000010";
      when "011001110110111" => color_data <= "000000000000";
      when "011001110111000" => color_data <= "000000000000";
      when "011001110111001" => color_data <= "000000000000";
      when "011001110111010" => color_data <= "000000000000";
      when "011001110111011" => color_data <= "000000000000";
      when "011001110111100" => color_data <= "000000000000";
      when "011001110111101" => color_data <= "000000000000";
      when "011001110111110" => color_data <= "000000000000";
      when "011001110111111" => color_data <= "000000000000";
      when "011001111000000" => color_data <= "000000000000";
      when "011001111000001" => color_data <= "000000000000";
      when "011001111000010" => color_data <= "000000000000";
      when "011001111000011" => color_data <= "000000000000";
      when "011001111000100" => color_data <= "000000000000";
      when "011001111000101" => color_data <= "000000000000";
      when "011001111000110" => color_data <= "000000000000";
      when "011001111000111" => color_data <= "000000000000";
      when "011001111001000" => color_data <= "000000000000";
      when "011001111001001" => color_data <= "000000000000";
      when "011001111001010" => color_data <= "000000000000";
      when "011001111001011" => color_data <= "000000000000";
      when "011001111001100" => color_data <= "000000000000";
      when "011001111001101" => color_data <= "000000000000";
      when "011001111001110" => color_data <= "000000000000";
      when "011001111001111" => color_data <= "000000000000";
      when "011001111010000" => color_data <= "000000000000";
      when "011001111010001" => color_data <= "000000000000";
      when "011001111010010" => color_data <= "000000000000";
      when "011001111010011" => color_data <= "000000000000";
      when "011001111010100" => color_data <= "000000000000";
      when "011001111010101" => color_data <= "000000000000";
      when "011001111010110" => color_data <= "000000000000";
      when "011001111010111" => color_data <= "000000000000";
      when "011001111011000" => color_data <= "000000000000";
      when "011001111011001" => color_data <= "000000000000";
      when "011001111011010" => color_data <= "000000000000";
      when "011001111011011" => color_data <= "000000000000";
      when "011001111011100" => color_data <= "000000000000";
      when "011001111011101" => color_data <= "000000000000";
      when "011001111011110" => color_data <= "000000000000";
      when "011001111011111" => color_data <= "000000000000";
      when "011001111100000" => color_data <= "000000000000";
      when "011001111100001" => color_data <= "000000000000";
      when "011001111100010" => color_data <= "000000000000";
      when "011001111100011" => color_data <= "000000000000";
      when "011010000000000" => color_data <= "000000000000";
      when "011010000000001" => color_data <= "000000000000";
      when "011010000000010" => color_data <= "000000000000";
      when "011010000000011" => color_data <= "000000000000";
      when "011010000000100" => color_data <= "000000000000";
      when "011010000000101" => color_data <= "000000000000";
      when "011010000000110" => color_data <= "000000000000";
      when "011010000000111" => color_data <= "000000000000";
      when "011010000001000" => color_data <= "000000000000";
      when "011010000001001" => color_data <= "000000000000";
      when "011010000001010" => color_data <= "000000000000";
      when "011010000001011" => color_data <= "000000000000";
      when "011010000001100" => color_data <= "000000000000";
      when "011010000001101" => color_data <= "000000000000";
      when "011010000001110" => color_data <= "000000000000";
      when "011010000001111" => color_data <= "000000000000";
      when "011010000010000" => color_data <= "000000000000";
      when "011010000010001" => color_data <= "000000000000";
      when "011010000010010" => color_data <= "000000000000";
      when "011010000010011" => color_data <= "000000000000";
      when "011010000010100" => color_data <= "000000000000";
      when "011010000010101" => color_data <= "000000000000";
      when "011010000010110" => color_data <= "000000000000";
      when "011010000010111" => color_data <= "000000000000";
      when "011010000011000" => color_data <= "000000000000";
      when "011010000011001" => color_data <= "000000000000";
      when "011010000011010" => color_data <= "000000000000";
      when "011010000011011" => color_data <= "000000000000";
      when "011010000011100" => color_data <= "000000000000";
      when "011010000011101" => color_data <= "000000000000";
      when "011010000011110" => color_data <= "000000000000";
      when "011010000011111" => color_data <= "000000000000";
      when "011010000100000" => color_data <= "000000000000";
      when "011010000100001" => color_data <= "000000000000";
      when "011010000100010" => color_data <= "000000000000";
      when "011010000100011" => color_data <= "000000000000";
      when "011010000100100" => color_data <= "000000000000";
      when "011010000100101" => color_data <= "000000000000";
      when "011010000100110" => color_data <= "000000000000";
      when "011010000100111" => color_data <= "000000000000";
      when "011010000101000" => color_data <= "000000000000";
      when "011010000101001" => color_data <= "000000000000";
      when "011010000101010" => color_data <= "000000000000";
      when "011010000101011" => color_data <= "000000000000";
      when "011010000101100" => color_data <= "000000000000";
      when "011010000101101" => color_data <= "000000000000";
      when "011010000101110" => color_data <= "011001010011";
      when "011010000101111" => color_data <= "111110110000";
      when "011010000110000" => color_data <= "111111000001";
      when "011010000110001" => color_data <= "111111000001";
      when "011010000110010" => color_data <= "111111000001";
      when "011010000110011" => color_data <= "111111000001";
      when "011010000110100" => color_data <= "111111000001";
      when "011010000110101" => color_data <= "111111000000";
      when "011010000110110" => color_data <= "101010000010";
      when "011010000110111" => color_data <= "000000000000";
      when "011010000111000" => color_data <= "000000000000";
      when "011010000111001" => color_data <= "000000000000";
      when "011010000111010" => color_data <= "000000000000";
      when "011010000111011" => color_data <= "000000000000";
      when "011010000111100" => color_data <= "000000000000";
      when "011010000111101" => color_data <= "000000000000";
      when "011010000111110" => color_data <= "000000000000";
      when "011010000111111" => color_data <= "000000000000";
      when "011010001000000" => color_data <= "000000000000";
      when "011010001000001" => color_data <= "000000000000";
      when "011010001000010" => color_data <= "000000000000";
      when "011010001000011" => color_data <= "000000000000";
      when "011010001000100" => color_data <= "000000000000";
      when "011010001000101" => color_data <= "000000000000";
      when "011010001000110" => color_data <= "000000000000";
      when "011010001000111" => color_data <= "000000000000";
      when "011010001001000" => color_data <= "000000000000";
      when "011010001001001" => color_data <= "000000000000";
      when "011010001001010" => color_data <= "000000000000";
      when "011010001001011" => color_data <= "000000000000";
      when "011010001001100" => color_data <= "000000000000";
      when "011010001001101" => color_data <= "000000000000";
      when "011010001001110" => color_data <= "000000000000";
      when "011010001001111" => color_data <= "000000000000";
      when "011010001010000" => color_data <= "000000000000";
      when "011010001010001" => color_data <= "000000000000";
      when "011010001010010" => color_data <= "000000000000";
      when "011010001010011" => color_data <= "000000000000";
      when "011010001010100" => color_data <= "000000000000";
      when "011010001010101" => color_data <= "000000000000";
      when "011010001010110" => color_data <= "000000000000";
      when "011010001010111" => color_data <= "000000000000";
      when "011010001011000" => color_data <= "000000000000";
      when "011010001011001" => color_data <= "000000000000";
      when "011010001011010" => color_data <= "000000000000";
      when "011010001011011" => color_data <= "000000000000";
      when "011010001011100" => color_data <= "000000000000";
      when "011010001011101" => color_data <= "000000000000";
      when "011010001011110" => color_data <= "000000000000";
      when "011010001011111" => color_data <= "000000000000";
      when "011010001100000" => color_data <= "000000000000";
      when "011010001100001" => color_data <= "000000000000";
      when "011010001100010" => color_data <= "000000000000";
      when "011010001100011" => color_data <= "000000000000";
      when "011010010000000" => color_data <= "000000000000";
      when "011010010000001" => color_data <= "000000000000";
      when "011010010000010" => color_data <= "000000000000";
      when "011010010000011" => color_data <= "000000000000";
      when "011010010000100" => color_data <= "000000000000";
      when "011010010000101" => color_data <= "000000000000";
      when "011010010000110" => color_data <= "000000000000";
      when "011010010000111" => color_data <= "000000000000";
      when "011010010001000" => color_data <= "000000000000";
      when "011010010001001" => color_data <= "000000000000";
      when "011010010001010" => color_data <= "000000000000";
      when "011010010001011" => color_data <= "000000000000";
      when "011010010001100" => color_data <= "000000000000";
      when "011010010001101" => color_data <= "000000000000";
      when "011010010001110" => color_data <= "000000000000";
      when "011010010001111" => color_data <= "000000000000";
      when "011010010010000" => color_data <= "000000000000";
      when "011010010010001" => color_data <= "000000000000";
      when "011010010010010" => color_data <= "000000000000";
      when "011010010010011" => color_data <= "000000000000";
      when "011010010010100" => color_data <= "000000000000";
      when "011010010010101" => color_data <= "000000000000";
      when "011010010010110" => color_data <= "000000000000";
      when "011010010010111" => color_data <= "000000000000";
      when "011010010011000" => color_data <= "000000000000";
      when "011010010011001" => color_data <= "000000000000";
      when "011010010011010" => color_data <= "000000000000";
      when "011010010011011" => color_data <= "000000000000";
      when "011010010011100" => color_data <= "000000000000";
      when "011010010011101" => color_data <= "000000000000";
      when "011010010011110" => color_data <= "000000000000";
      when "011010010011111" => color_data <= "000000000000";
      when "011010010100000" => color_data <= "000000000000";
      when "011010010100001" => color_data <= "000000000000";
      when "011010010100010" => color_data <= "000000000000";
      when "011010010100011" => color_data <= "000000000000";
      when "011010010100100" => color_data <= "000000000000";
      when "011010010100101" => color_data <= "000000000000";
      when "011010010100110" => color_data <= "000000000000";
      when "011010010100111" => color_data <= "000000000000";
      when "011010010101000" => color_data <= "000000000000";
      when "011010010101001" => color_data <= "000000000000";
      when "011010010101010" => color_data <= "000000000000";
      when "011010010101011" => color_data <= "000000000000";
      when "011010010101100" => color_data <= "000000000000";
      when "011010010101101" => color_data <= "000000000000";
      when "011010010101110" => color_data <= "011101100011";
      when "011010010101111" => color_data <= "111110110000";
      when "011010010110000" => color_data <= "111111000001";
      when "011010010110001" => color_data <= "111111000001";
      when "011010010110010" => color_data <= "111111000001";
      when "011010010110011" => color_data <= "111111000001";
      when "011010010110100" => color_data <= "111111000001";
      when "011010010110101" => color_data <= "111111000000";
      when "011010010110110" => color_data <= "101110010001";
      when "011010010110111" => color_data <= "000000000000";
      when "011010010111000" => color_data <= "000000000000";
      when "011010010111001" => color_data <= "000000000000";
      when "011010010111010" => color_data <= "000000000000";
      when "011010010111011" => color_data <= "000000000000";
      when "011010010111100" => color_data <= "000000000000";
      when "011010010111101" => color_data <= "000000000000";
      when "011010010111110" => color_data <= "000000000000";
      when "011010010111111" => color_data <= "000000000000";
      when "011010011000000" => color_data <= "000000000000";
      when "011010011000001" => color_data <= "000000000000";
      when "011010011000010" => color_data <= "000000000000";
      when "011010011000011" => color_data <= "000000000000";
      when "011010011000100" => color_data <= "000000000000";
      when "011010011000101" => color_data <= "000000000000";
      when "011010011000110" => color_data <= "000000000000";
      when "011010011000111" => color_data <= "000000000000";
      when "011010011001000" => color_data <= "000000000000";
      when "011010011001001" => color_data <= "000000000000";
      when "011010011001010" => color_data <= "000000000000";
      when "011010011001011" => color_data <= "000000000000";
      when "011010011001100" => color_data <= "000000000000";
      when "011010011001101" => color_data <= "000000000000";
      when "011010011001110" => color_data <= "000000000000";
      when "011010011001111" => color_data <= "000000000000";
      when "011010011010000" => color_data <= "000000000000";
      when "011010011010001" => color_data <= "000000000000";
      when "011010011010010" => color_data <= "000000000000";
      when "011010011010011" => color_data <= "000000000000";
      when "011010011010100" => color_data <= "000000000000";
      when "011010011010101" => color_data <= "000000000000";
      when "011010011010110" => color_data <= "000000000000";
      when "011010011010111" => color_data <= "000000000000";
      when "011010011011000" => color_data <= "000000000000";
      when "011010011011001" => color_data <= "000000000000";
      when "011010011011010" => color_data <= "000000000000";
      when "011010011011011" => color_data <= "000000000000";
      when "011010011011100" => color_data <= "000000000000";
      when "011010011011101" => color_data <= "000000000000";
      when "011010011011110" => color_data <= "000000000000";
      when "011010011011111" => color_data <= "000000000000";
      when "011010011100000" => color_data <= "000000000000";
      when "011010011100001" => color_data <= "000000000000";
      when "011010011100010" => color_data <= "000000000000";
      when "011010011100011" => color_data <= "000000000000";
      when "011010100000000" => color_data <= "000000000000";
      when "011010100000001" => color_data <= "000000000000";
      when "011010100000010" => color_data <= "000000000000";
      when "011010100000011" => color_data <= "000000000000";
      when "011010100000100" => color_data <= "000000000000";
      when "011010100000101" => color_data <= "000000000000";
      when "011010100000110" => color_data <= "000000000000";
      when "011010100000111" => color_data <= "000000000000";
      when "011010100001000" => color_data <= "000000000000";
      when "011010100001001" => color_data <= "000000000000";
      when "011010100001010" => color_data <= "000000000000";
      when "011010100001011" => color_data <= "000000000000";
      when "011010100001100" => color_data <= "000000000000";
      when "011010100001101" => color_data <= "000000000000";
      when "011010100001110" => color_data <= "000000000000";
      when "011010100001111" => color_data <= "000000000000";
      when "011010100010000" => color_data <= "000000000000";
      when "011010100010001" => color_data <= "000000000000";
      when "011010100010010" => color_data <= "000000000000";
      when "011010100010011" => color_data <= "000000000000";
      when "011010100010100" => color_data <= "000000000000";
      when "011010100010101" => color_data <= "000000000000";
      when "011010100010110" => color_data <= "000000000000";
      when "011010100010111" => color_data <= "000000000000";
      when "011010100011000" => color_data <= "000000000000";
      when "011010100011001" => color_data <= "000000000000";
      when "011010100011010" => color_data <= "000000000000";
      when "011010100011011" => color_data <= "000000000000";
      when "011010100011100" => color_data <= "000000000000";
      when "011010100011101" => color_data <= "000000000000";
      when "011010100011110" => color_data <= "000000000000";
      when "011010100011111" => color_data <= "000000000000";
      when "011010100100000" => color_data <= "000000000000";
      when "011010100100001" => color_data <= "000000000000";
      when "011010100100010" => color_data <= "000000000000";
      when "011010100100011" => color_data <= "000000000000";
      when "011010100100100" => color_data <= "000000000000";
      when "011010100100101" => color_data <= "000000000000";
      when "011010100100110" => color_data <= "000000000000";
      when "011010100100111" => color_data <= "000000000000";
      when "011010100101000" => color_data <= "000000000000";
      when "011010100101001" => color_data <= "000000000000";
      when "011010100101010" => color_data <= "000000000000";
      when "011010100101011" => color_data <= "000000000000";
      when "011010100101100" => color_data <= "000000000000";
      when "011010100101101" => color_data <= "000000000000";
      when "011010100101110" => color_data <= "100001110010";
      when "011010100101111" => color_data <= "111110110000";
      when "011010100110000" => color_data <= "111111000001";
      when "011010100110001" => color_data <= "111111000001";
      when "011010100110010" => color_data <= "111111000001";
      when "011010100110011" => color_data <= "111111000001";
      when "011010100110100" => color_data <= "111111000001";
      when "011010100110101" => color_data <= "111111000000";
      when "011010100110110" => color_data <= "110010010000";
      when "011010100110111" => color_data <= "000000000000";
      when "011010100111000" => color_data <= "000000000000";
      when "011010100111001" => color_data <= "000000000000";
      when "011010100111010" => color_data <= "000000000000";
      when "011010100111011" => color_data <= "000000000000";
      when "011010100111100" => color_data <= "000000000000";
      when "011010100111101" => color_data <= "000000000000";
      when "011010100111110" => color_data <= "000000000000";
      when "011010100111111" => color_data <= "000000000000";
      when "011010101000000" => color_data <= "000000000000";
      when "011010101000001" => color_data <= "000000000000";
      when "011010101000010" => color_data <= "000000000000";
      when "011010101000011" => color_data <= "000000000000";
      when "011010101000100" => color_data <= "000000000000";
      when "011010101000101" => color_data <= "000000000000";
      when "011010101000110" => color_data <= "000000000000";
      when "011010101000111" => color_data <= "000000000000";
      when "011010101001000" => color_data <= "000000000000";
      when "011010101001001" => color_data <= "000000000000";
      when "011010101001010" => color_data <= "000000000000";
      when "011010101001011" => color_data <= "000000000000";
      when "011010101001100" => color_data <= "000000000000";
      when "011010101001101" => color_data <= "000000000000";
      when "011010101001110" => color_data <= "000000000000";
      when "011010101001111" => color_data <= "000000000000";
      when "011010101010000" => color_data <= "000000000000";
      when "011010101010001" => color_data <= "000000000000";
      when "011010101010010" => color_data <= "000000000000";
      when "011010101010011" => color_data <= "000000000000";
      when "011010101010100" => color_data <= "000000000000";
      when "011010101010101" => color_data <= "000000000000";
      when "011010101010110" => color_data <= "000000000000";
      when "011010101010111" => color_data <= "000000000000";
      when "011010101011000" => color_data <= "000000000000";
      when "011010101011001" => color_data <= "000000000000";
      when "011010101011010" => color_data <= "000000000000";
      when "011010101011011" => color_data <= "000000000000";
      when "011010101011100" => color_data <= "000000000000";
      when "011010101011101" => color_data <= "000000000000";
      when "011010101011110" => color_data <= "000000000000";
      when "011010101011111" => color_data <= "000000000000";
      when "011010101100000" => color_data <= "000000000000";
      when "011010101100001" => color_data <= "000000000000";
      when "011010101100010" => color_data <= "000000000000";
      when "011010101100011" => color_data <= "000000000000";
      when "011010110000000" => color_data <= "000000000000";
      when "011010110000001" => color_data <= "000000000000";
      when "011010110000010" => color_data <= "000000000000";
      when "011010110000011" => color_data <= "000000000000";
      when "011010110000100" => color_data <= "000000000000";
      when "011010110000101" => color_data <= "000000000000";
      when "011010110000110" => color_data <= "000000000000";
      when "011010110000111" => color_data <= "000000000000";
      when "011010110001000" => color_data <= "000000000000";
      when "011010110001001" => color_data <= "000000000000";
      when "011010110001010" => color_data <= "000000000000";
      when "011010110001011" => color_data <= "000000000000";
      when "011010110001100" => color_data <= "000000000000";
      when "011010110001101" => color_data <= "000000000000";
      when "011010110001110" => color_data <= "000000000000";
      when "011010110001111" => color_data <= "000000000000";
      when "011010110010000" => color_data <= "000000000000";
      when "011010110010001" => color_data <= "000000000000";
      when "011010110010010" => color_data <= "000000000000";
      when "011010110010011" => color_data <= "000000000000";
      when "011010110010100" => color_data <= "000000000000";
      when "011010110010101" => color_data <= "000000000000";
      when "011010110010110" => color_data <= "000000000000";
      when "011010110010111" => color_data <= "000000000000";
      when "011010110011000" => color_data <= "000000000000";
      when "011010110011001" => color_data <= "000000000000";
      when "011010110011010" => color_data <= "000000000000";
      when "011010110011011" => color_data <= "000000000000";
      when "011010110011100" => color_data <= "000000000000";
      when "011010110011101" => color_data <= "000000000000";
      when "011010110011110" => color_data <= "000000000000";
      when "011010110011111" => color_data <= "000000000000";
      when "011010110100000" => color_data <= "000000000000";
      when "011010110100001" => color_data <= "000000000000";
      when "011010110100010" => color_data <= "000000000000";
      when "011010110100011" => color_data <= "000000000000";
      when "011010110100100" => color_data <= "000000000000";
      when "011010110100101" => color_data <= "000000000000";
      when "011010110100110" => color_data <= "000000000000";
      when "011010110100111" => color_data <= "000000000000";
      when "011010110101000" => color_data <= "000000000000";
      when "011010110101001" => color_data <= "000000000000";
      when "011010110101010" => color_data <= "000000000000";
      when "011010110101011" => color_data <= "000000000000";
      when "011010110101100" => color_data <= "000000000000";
      when "011010110101101" => color_data <= "000000000000";
      when "011010110101110" => color_data <= "101010000010";
      when "011010110101111" => color_data <= "111111000000";
      when "011010110110000" => color_data <= "111111000001";
      when "011010110110001" => color_data <= "111111000001";
      when "011010110110010" => color_data <= "111111000000";
      when "011010110110011" => color_data <= "111111000000";
      when "011010110110100" => color_data <= "111111000000";
      when "011010110110101" => color_data <= "111111000001";
      when "011010110110110" => color_data <= "111111000000";
      when "011010110110111" => color_data <= "000100010001";
      when "011010110111000" => color_data <= "000000000000";
      when "011010110111001" => color_data <= "000000000000";
      when "011010110111010" => color_data <= "000000000000";
      when "011010110111011" => color_data <= "000000000000";
      when "011010110111100" => color_data <= "000000000000";
      when "011010110111101" => color_data <= "000000000000";
      when "011010110111110" => color_data <= "000000000000";
      when "011010110111111" => color_data <= "000000000000";
      when "011010111000000" => color_data <= "000000000000";
      when "011010111000001" => color_data <= "000000000000";
      when "011010111000010" => color_data <= "000000000000";
      when "011010111000011" => color_data <= "000000000000";
      when "011010111000100" => color_data <= "000000000000";
      when "011010111000101" => color_data <= "000000000000";
      when "011010111000110" => color_data <= "000000000000";
      when "011010111000111" => color_data <= "000000000000";
      when "011010111001000" => color_data <= "000000000000";
      when "011010111001001" => color_data <= "000000000000";
      when "011010111001010" => color_data <= "000000000000";
      when "011010111001011" => color_data <= "000000000000";
      when "011010111001100" => color_data <= "000000000000";
      when "011010111001101" => color_data <= "000000000000";
      when "011010111001110" => color_data <= "000000000000";
      when "011010111001111" => color_data <= "000000000000";
      when "011010111010000" => color_data <= "000000000000";
      when "011010111010001" => color_data <= "000000000000";
      when "011010111010010" => color_data <= "000000000000";
      when "011010111010011" => color_data <= "000000000000";
      when "011010111010100" => color_data <= "000000000000";
      when "011010111010101" => color_data <= "000000000000";
      when "011010111010110" => color_data <= "000000000000";
      when "011010111010111" => color_data <= "000000000000";
      when "011010111011000" => color_data <= "000000000000";
      when "011010111011001" => color_data <= "000000000000";
      when "011010111011010" => color_data <= "000000000000";
      when "011010111011011" => color_data <= "000000000000";
      when "011010111011100" => color_data <= "000000000000";
      when "011010111011101" => color_data <= "000000000000";
      when "011010111011110" => color_data <= "000000000000";
      when "011010111011111" => color_data <= "000000000000";
      when "011010111100000" => color_data <= "000000000000";
      when "011010111100001" => color_data <= "000000000000";
      when "011010111100010" => color_data <= "000000000000";
      when "011010111100011" => color_data <= "000000000000";
      when "011011000000000" => color_data <= "000000000000";
      when "011011000000001" => color_data <= "000000000000";
      when "011011000000010" => color_data <= "000000000000";
      when "011011000000011" => color_data <= "000000000000";
      when "011011000000100" => color_data <= "000000000000";
      when "011011000000101" => color_data <= "000000000000";
      when "011011000000110" => color_data <= "000000000000";
      when "011011000000111" => color_data <= "000000000000";
      when "011011000001000" => color_data <= "000000000000";
      when "011011000001001" => color_data <= "000000000000";
      when "011011000001010" => color_data <= "000000000000";
      when "011011000001011" => color_data <= "000000000000";
      when "011011000001100" => color_data <= "000000000000";
      when "011011000001101" => color_data <= "000000000000";
      when "011011000001110" => color_data <= "000000000000";
      when "011011000001111" => color_data <= "000000000000";
      when "011011000010000" => color_data <= "000000000000";
      when "011011000010001" => color_data <= "000000000000";
      when "011011000010010" => color_data <= "000000000000";
      when "011011000010011" => color_data <= "000000000000";
      when "011011000010100" => color_data <= "000000000000";
      when "011011000010101" => color_data <= "000000000000";
      when "011011000010110" => color_data <= "000000000000";
      when "011011000010111" => color_data <= "000000000000";
      when "011011000011000" => color_data <= "000000000000";
      when "011011000011001" => color_data <= "000000000000";
      when "011011000011010" => color_data <= "000000000000";
      when "011011000011011" => color_data <= "000000000000";
      when "011011000011100" => color_data <= "000000000000";
      when "011011000011101" => color_data <= "000000000000";
      when "011011000011110" => color_data <= "000000000000";
      when "011011000011111" => color_data <= "000000000000";
      when "011011000100000" => color_data <= "000000000000";
      when "011011000100001" => color_data <= "000000000000";
      when "011011000100010" => color_data <= "000000000000";
      when "011011000100011" => color_data <= "000000000000";
      when "011011000100100" => color_data <= "000000000000";
      when "011011000100101" => color_data <= "000000000000";
      when "011011000100110" => color_data <= "000000000000";
      when "011011000100111" => color_data <= "000000000000";
      when "011011000101000" => color_data <= "000000000000";
      when "011011000101001" => color_data <= "000000000000";
      when "011011000101010" => color_data <= "000000000000";
      when "011011000101011" => color_data <= "000000000000";
      when "011011000101100" => color_data <= "000000000000";
      when "011011000101101" => color_data <= "000000000000";
      when "011011000101110" => color_data <= "101110010001";
      when "011011000101111" => color_data <= "111111000000";
      when "011011000110000" => color_data <= "111111000001";
      when "011011000110001" => color_data <= "111111000000";
      when "011011000110010" => color_data <= "111111000011";
      when "011011000110011" => color_data <= "111111010110";
      when "011011000110100" => color_data <= "111111000010";
      when "011011000110101" => color_data <= "111111000000";
      when "011011000110110" => color_data <= "111110110000";
      when "011011000110111" => color_data <= "001000100010";
      when "011011000111000" => color_data <= "000000000000";
      when "011011000111001" => color_data <= "000000000000";
      when "011011000111010" => color_data <= "000000000000";
      when "011011000111011" => color_data <= "000000000000";
      when "011011000111100" => color_data <= "000000000000";
      when "011011000111101" => color_data <= "000000000000";
      when "011011000111110" => color_data <= "000000000000";
      when "011011000111111" => color_data <= "000000000000";
      when "011011001000000" => color_data <= "000000000000";
      when "011011001000001" => color_data <= "000000000000";
      when "011011001000010" => color_data <= "000000000000";
      when "011011001000011" => color_data <= "000000000000";
      when "011011001000100" => color_data <= "000000000000";
      when "011011001000101" => color_data <= "000000000000";
      when "011011001000110" => color_data <= "000000000000";
      when "011011001000111" => color_data <= "000000000000";
      when "011011001001000" => color_data <= "000000000000";
      when "011011001001001" => color_data <= "000000000000";
      when "011011001001010" => color_data <= "000000000000";
      when "011011001001011" => color_data <= "000000000000";
      when "011011001001100" => color_data <= "000000000000";
      when "011011001001101" => color_data <= "000000000000";
      when "011011001001110" => color_data <= "000000000000";
      when "011011001001111" => color_data <= "000000000000";
      when "011011001010000" => color_data <= "000000000000";
      when "011011001010001" => color_data <= "000000000000";
      when "011011001010010" => color_data <= "000000000000";
      when "011011001010011" => color_data <= "000000000000";
      when "011011001010100" => color_data <= "000000000000";
      when "011011001010101" => color_data <= "000000000000";
      when "011011001010110" => color_data <= "000000000000";
      when "011011001010111" => color_data <= "000000000000";
      when "011011001011000" => color_data <= "000000000000";
      when "011011001011001" => color_data <= "000000000000";
      when "011011001011010" => color_data <= "000000000000";
      when "011011001011011" => color_data <= "000000000000";
      when "011011001011100" => color_data <= "000000000000";
      when "011011001011101" => color_data <= "000000000000";
      when "011011001011110" => color_data <= "000000000000";
      when "011011001011111" => color_data <= "000000000000";
      when "011011001100000" => color_data <= "000000000000";
      when "011011001100001" => color_data <= "000000000000";
      when "011011001100010" => color_data <= "000000000000";
      when "011011001100011" => color_data <= "000000000000";
      when "011011010000000" => color_data <= "000000000000";
      when "011011010000001" => color_data <= "000000000000";
      when "011011010000010" => color_data <= "000000000000";
      when "011011010000011" => color_data <= "000000000000";
      when "011011010000100" => color_data <= "000000000000";
      when "011011010000101" => color_data <= "000000000000";
      when "011011010000110" => color_data <= "000000000000";
      when "011011010000111" => color_data <= "000000000000";
      when "011011010001000" => color_data <= "000000000000";
      when "011011010001001" => color_data <= "000000000000";
      when "011011010001010" => color_data <= "000000000000";
      when "011011010001011" => color_data <= "000000000000";
      when "011011010001100" => color_data <= "000000000000";
      when "011011010001101" => color_data <= "000000000000";
      when "011011010001110" => color_data <= "000000000000";
      when "011011010001111" => color_data <= "000000000000";
      when "011011010010000" => color_data <= "000000000000";
      when "011011010010001" => color_data <= "000000000000";
      when "011011010010010" => color_data <= "000000000000";
      when "011011010010011" => color_data <= "000000000000";
      when "011011010010100" => color_data <= "000000000000";
      when "011011010010101" => color_data <= "000000000000";
      when "011011010010110" => color_data <= "000000000000";
      when "011011010010111" => color_data <= "000000000000";
      when "011011010011000" => color_data <= "000000000000";
      when "011011010011001" => color_data <= "000000000000";
      when "011011010011010" => color_data <= "000000000000";
      when "011011010011011" => color_data <= "000000000000";
      when "011011010011100" => color_data <= "000000000000";
      when "011011010011101" => color_data <= "000000000000";
      when "011011010011110" => color_data <= "000000000000";
      when "011011010011111" => color_data <= "000000000000";
      when "011011010100000" => color_data <= "000000000000";
      when "011011010100001" => color_data <= "000000000000";
      when "011011010100010" => color_data <= "000000000000";
      when "011011010100011" => color_data <= "000000000000";
      when "011011010100100" => color_data <= "000000000000";
      when "011011010100101" => color_data <= "000000000000";
      when "011011010100110" => color_data <= "000000000000";
      when "011011010100111" => color_data <= "000000000000";
      when "011011010101000" => color_data <= "000000000000";
      when "011011010101001" => color_data <= "000000000000";
      when "011011010101010" => color_data <= "000000000000";
      when "011011010101011" => color_data <= "000000000000";
      when "011011010101100" => color_data <= "000000000000";
      when "011011010101101" => color_data <= "000000000000";
      when "011011010101110" => color_data <= "110110100000";
      when "011011010101111" => color_data <= "111111000000";
      when "011011010110000" => color_data <= "111111000001";
      when "011011010110001" => color_data <= "111111000000";
      when "011011010110010" => color_data <= "111111000011";
      when "011011010110011" => color_data <= "111111101001";
      when "011011010110100" => color_data <= "111111010100";
      when "011011010110101" => color_data <= "111111000000";
      when "011011010110110" => color_data <= "111110110000";
      when "011011010110111" => color_data <= "001100110010";
      when "011011010111000" => color_data <= "000000000000";
      when "011011010111001" => color_data <= "000000000000";
      when "011011010111010" => color_data <= "000000000000";
      when "011011010111011" => color_data <= "000000000000";
      when "011011010111100" => color_data <= "000000000000";
      when "011011010111101" => color_data <= "000000000000";
      when "011011010111110" => color_data <= "000000000000";
      when "011011010111111" => color_data <= "000000000000";
      when "011011011000000" => color_data <= "000000000000";
      when "011011011000001" => color_data <= "000000000000";
      when "011011011000010" => color_data <= "000000000000";
      when "011011011000011" => color_data <= "000000000000";
      when "011011011000100" => color_data <= "000000000000";
      when "011011011000101" => color_data <= "000000000000";
      when "011011011000110" => color_data <= "000000000000";
      when "011011011000111" => color_data <= "000000000000";
      when "011011011001000" => color_data <= "000000000000";
      when "011011011001001" => color_data <= "000000000000";
      when "011011011001010" => color_data <= "000000000000";
      when "011011011001011" => color_data <= "000000000000";
      when "011011011001100" => color_data <= "000000000000";
      when "011011011001101" => color_data <= "000000000000";
      when "011011011001110" => color_data <= "000000000000";
      when "011011011001111" => color_data <= "000000000000";
      when "011011011010000" => color_data <= "000000000000";
      when "011011011010001" => color_data <= "000000000000";
      when "011011011010010" => color_data <= "000000000000";
      when "011011011010011" => color_data <= "000000000000";
      when "011011011010100" => color_data <= "000000000000";
      when "011011011010101" => color_data <= "000000000000";
      when "011011011010110" => color_data <= "000000000000";
      when "011011011010111" => color_data <= "000000000000";
      when "011011011011000" => color_data <= "000000000000";
      when "011011011011001" => color_data <= "000000000000";
      when "011011011011010" => color_data <= "000000000000";
      when "011011011011011" => color_data <= "000000000000";
      when "011011011011100" => color_data <= "000000000000";
      when "011011011011101" => color_data <= "000000000000";
      when "011011011011110" => color_data <= "000000000000";
      when "011011011011111" => color_data <= "000000000000";
      when "011011011100000" => color_data <= "000000000000";
      when "011011011100001" => color_data <= "000000000000";
      when "011011011100010" => color_data <= "000000000000";
      when "011011011100011" => color_data <= "000000000000";
      when "011011100000000" => color_data <= "000000000000";
      when "011011100000001" => color_data <= "000000000000";
      when "011011100000010" => color_data <= "000000000000";
      when "011011100000011" => color_data <= "000000000000";
      when "011011100000100" => color_data <= "000000000000";
      when "011011100000101" => color_data <= "000000000000";
      when "011011100000110" => color_data <= "000000000000";
      when "011011100000111" => color_data <= "000000000000";
      when "011011100001000" => color_data <= "000000000000";
      when "011011100001001" => color_data <= "000000000000";
      when "011011100001010" => color_data <= "000000000000";
      when "011011100001011" => color_data <= "000000000000";
      when "011011100001100" => color_data <= "000000000000";
      when "011011100001101" => color_data <= "000000000000";
      when "011011100001110" => color_data <= "000000000000";
      when "011011100001111" => color_data <= "000000000000";
      when "011011100010000" => color_data <= "000000000000";
      when "011011100010001" => color_data <= "000000000000";
      when "011011100010010" => color_data <= "000000000000";
      when "011011100010011" => color_data <= "000000000000";
      when "011011100010100" => color_data <= "000000000000";
      when "011011100010101" => color_data <= "000000000000";
      when "011011100010110" => color_data <= "000000000000";
      when "011011100010111" => color_data <= "000000000000";
      when "011011100011000" => color_data <= "000000000000";
      when "011011100011001" => color_data <= "000000000000";
      when "011011100011010" => color_data <= "000000000000";
      when "011011100011011" => color_data <= "000000000000";
      when "011011100011100" => color_data <= "000000000000";
      when "011011100011101" => color_data <= "000000000000";
      when "011011100011110" => color_data <= "000000000000";
      when "011011100011111" => color_data <= "000000000000";
      when "011011100100000" => color_data <= "000000000000";
      when "011011100100001" => color_data <= "000000000000";
      when "011011100100010" => color_data <= "000000000000";
      when "011011100100011" => color_data <= "000000000000";
      when "011011100100100" => color_data <= "000000000000";
      when "011011100100101" => color_data <= "000000000000";
      when "011011100100110" => color_data <= "000000000000";
      when "011011100100111" => color_data <= "000000000000";
      when "011011100101000" => color_data <= "000000000000";
      when "011011100101001" => color_data <= "000000000000";
      when "011011100101010" => color_data <= "000000000000";
      when "011011100101011" => color_data <= "000000000000";
      when "011011100101100" => color_data <= "001000100001";
      when "011011100101101" => color_data <= "010101010011";
      when "011011100101110" => color_data <= "110110100000";
      when "011011100101111" => color_data <= "111111000001";
      when "011011100110000" => color_data <= "111111000001";
      when "011011100110001" => color_data <= "111111000000";
      when "011011100110010" => color_data <= "111111010100";
      when "011011100110011" => color_data <= "111111101010";
      when "011011100110100" => color_data <= "111111010100";
      when "011011100110101" => color_data <= "111111000000";
      when "011011100110110" => color_data <= "111110110000";
      when "011011100110111" => color_data <= "100001110010";
      when "011011100111000" => color_data <= "001000100001";
      when "011011100111001" => color_data <= "000000000000";
      when "011011100111010" => color_data <= "000000000000";
      when "011011100111011" => color_data <= "000000000000";
      when "011011100111100" => color_data <= "000000000000";
      when "011011100111101" => color_data <= "000000000000";
      when "011011100111110" => color_data <= "000000000000";
      when "011011100111111" => color_data <= "000000000000";
      when "011011101000000" => color_data <= "000000000000";
      when "011011101000001" => color_data <= "000000000000";
      when "011011101000010" => color_data <= "000000000000";
      when "011011101000011" => color_data <= "000000000000";
      when "011011101000100" => color_data <= "000000000000";
      when "011011101000101" => color_data <= "000000000000";
      when "011011101000110" => color_data <= "000000000000";
      when "011011101000111" => color_data <= "000000000000";
      when "011011101001000" => color_data <= "000000000000";
      when "011011101001001" => color_data <= "000000000000";
      when "011011101001010" => color_data <= "000000000000";
      when "011011101001011" => color_data <= "000000000000";
      when "011011101001100" => color_data <= "000000000000";
      when "011011101001101" => color_data <= "000000000000";
      when "011011101001110" => color_data <= "000000000000";
      when "011011101001111" => color_data <= "000000000000";
      when "011011101010000" => color_data <= "000000000000";
      when "011011101010001" => color_data <= "000000000000";
      when "011011101010010" => color_data <= "000000000000";
      when "011011101010011" => color_data <= "000000000000";
      when "011011101010100" => color_data <= "000000000000";
      when "011011101010101" => color_data <= "000000000000";
      when "011011101010110" => color_data <= "000000000000";
      when "011011101010111" => color_data <= "000000000000";
      when "011011101011000" => color_data <= "000000000000";
      when "011011101011001" => color_data <= "000000000000";
      when "011011101011010" => color_data <= "000000000000";
      when "011011101011011" => color_data <= "000000000000";
      when "011011101011100" => color_data <= "000000000000";
      when "011011101011101" => color_data <= "000000000000";
      when "011011101011110" => color_data <= "000000000000";
      when "011011101011111" => color_data <= "000000000000";
      when "011011101100000" => color_data <= "000000000000";
      when "011011101100001" => color_data <= "000000000000";
      when "011011101100010" => color_data <= "000000000000";
      when "011011101100011" => color_data <= "000000000000";
      when "011011110000000" => color_data <= "000000000000";
      when "011011110000001" => color_data <= "000000000000";
      when "011011110000010" => color_data <= "000000000000";
      when "011011110000011" => color_data <= "000000000000";
      when "011011110000100" => color_data <= "000000000000";
      when "011011110000101" => color_data <= "000000000000";
      when "011011110000110" => color_data <= "000000000000";
      when "011011110000111" => color_data <= "000000000000";
      when "011011110001000" => color_data <= "000000000000";
      when "011011110001001" => color_data <= "000000000000";
      when "011011110001010" => color_data <= "000000000000";
      when "011011110001011" => color_data <= "000000000000";
      when "011011110001100" => color_data <= "000000000000";
      when "011011110001101" => color_data <= "000000000000";
      when "011011110001110" => color_data <= "000000000000";
      when "011011110001111" => color_data <= "000000000000";
      when "011011110010000" => color_data <= "000000000000";
      when "011011110010001" => color_data <= "000000000000";
      when "011011110010010" => color_data <= "000000000000";
      when "011011110010011" => color_data <= "000000000000";
      when "011011110010100" => color_data <= "000000000000";
      when "011011110010101" => color_data <= "000000000000";
      when "011011110010110" => color_data <= "000000000000";
      when "011011110010111" => color_data <= "000000000000";
      when "011011110011000" => color_data <= "000000000000";
      when "011011110011001" => color_data <= "000000000000";
      when "011011110011010" => color_data <= "000000000000";
      when "011011110011011" => color_data <= "000000000000";
      when "011011110011100" => color_data <= "000000000000";
      when "011011110011101" => color_data <= "000000000000";
      when "011011110011110" => color_data <= "000000000000";
      when "011011110011111" => color_data <= "000000000000";
      when "011011110100000" => color_data <= "000000000000";
      when "011011110100001" => color_data <= "000000000000";
      when "011011110100010" => color_data <= "000000000000";
      when "011011110100011" => color_data <= "000000000000";
      when "011011110100100" => color_data <= "000000000000";
      when "011011110100101" => color_data <= "000000000000";
      when "011011110100110" => color_data <= "000000000000";
      when "011011110100111" => color_data <= "000000000000";
      when "011011110101000" => color_data <= "000000000000";
      when "011011110101001" => color_data <= "000000000000";
      when "011011110101010" => color_data <= "000000000000";
      when "011011110101011" => color_data <= "000000000000";
      when "011011110101100" => color_data <= "011101100011";
      when "011011110101101" => color_data <= "111110110000";
      when "011011110101110" => color_data <= "111111000001";
      when "011011110101111" => color_data <= "111111000001";
      when "011011110110000" => color_data <= "111111000001";
      when "011011110110001" => color_data <= "111111000000";
      when "011011110110010" => color_data <= "111111000010";
      when "011011110110011" => color_data <= "111111010100";
      when "011011110110100" => color_data <= "111111000010";
      when "011011110110101" => color_data <= "111111000001";
      when "011011110110110" => color_data <= "111111000001";
      when "011011110110111" => color_data <= "111110110000";
      when "011011110111000" => color_data <= "100001110010";
      when "011011110111001" => color_data <= "000000000000";
      when "011011110111010" => color_data <= "000000000000";
      when "011011110111011" => color_data <= "000000000000";
      when "011011110111100" => color_data <= "000000000000";
      when "011011110111101" => color_data <= "000000000000";
      when "011011110111110" => color_data <= "000000000000";
      when "011011110111111" => color_data <= "000000000000";
      when "011011111000000" => color_data <= "000000000000";
      when "011011111000001" => color_data <= "000000000000";
      when "011011111000010" => color_data <= "000000000000";
      when "011011111000011" => color_data <= "000000000000";
      when "011011111000100" => color_data <= "000000000000";
      when "011011111000101" => color_data <= "000000000000";
      when "011011111000110" => color_data <= "000000000000";
      when "011011111000111" => color_data <= "000000000000";
      when "011011111001000" => color_data <= "000000000000";
      when "011011111001001" => color_data <= "000000000000";
      when "011011111001010" => color_data <= "000000000000";
      when "011011111001011" => color_data <= "000000000000";
      when "011011111001100" => color_data <= "000000000000";
      when "011011111001101" => color_data <= "000000000000";
      when "011011111001110" => color_data <= "000000000000";
      when "011011111001111" => color_data <= "000000000000";
      when "011011111010000" => color_data <= "000000000000";
      when "011011111010001" => color_data <= "000000000000";
      when "011011111010010" => color_data <= "000000000000";
      when "011011111010011" => color_data <= "000000000000";
      when "011011111010100" => color_data <= "000000000000";
      when "011011111010101" => color_data <= "000000000000";
      when "011011111010110" => color_data <= "000000000000";
      when "011011111010111" => color_data <= "000000000000";
      when "011011111011000" => color_data <= "000000000000";
      when "011011111011001" => color_data <= "000000000000";
      when "011011111011010" => color_data <= "000000000000";
      when "011011111011011" => color_data <= "000000000000";
      when "011011111011100" => color_data <= "000000000000";
      when "011011111011101" => color_data <= "000000000000";
      when "011011111011110" => color_data <= "000000000000";
      when "011011111011111" => color_data <= "000000000000";
      when "011011111100000" => color_data <= "000000000000";
      when "011011111100001" => color_data <= "000000000000";
      when "011011111100010" => color_data <= "000000000000";
      when "011011111100011" => color_data <= "000000000000";
      when "011100000000000" => color_data <= "000000000000";
      when "011100000000001" => color_data <= "000000000000";
      when "011100000000010" => color_data <= "000000000000";
      when "011100000000011" => color_data <= "000000000000";
      when "011100000000100" => color_data <= "000000000000";
      when "011100000000101" => color_data <= "000000000000";
      when "011100000000110" => color_data <= "000000000000";
      when "011100000000111" => color_data <= "000000000000";
      when "011100000001000" => color_data <= "000000000000";
      when "011100000001001" => color_data <= "000000000000";
      when "011100000001010" => color_data <= "000000000000";
      when "011100000001011" => color_data <= "000000000000";
      when "011100000001100" => color_data <= "000000000000";
      when "011100000001101" => color_data <= "000000000000";
      when "011100000001110" => color_data <= "000000000000";
      when "011100000001111" => color_data <= "000000000000";
      when "011100000010000" => color_data <= "000000000000";
      when "011100000010001" => color_data <= "000000000000";
      when "011100000010010" => color_data <= "000000000000";
      when "011100000010011" => color_data <= "000000000000";
      when "011100000010100" => color_data <= "000000000000";
      when "011100000010101" => color_data <= "000000000000";
      when "011100000010110" => color_data <= "000000000000";
      when "011100000010111" => color_data <= "000000000000";
      when "011100000011000" => color_data <= "000000000000";
      when "011100000011001" => color_data <= "000000000000";
      when "011100000011010" => color_data <= "000000000000";
      when "011100000011011" => color_data <= "000000000000";
      when "011100000011100" => color_data <= "000000000000";
      when "011100000011101" => color_data <= "000000000000";
      when "011100000011110" => color_data <= "000000000000";
      when "011100000011111" => color_data <= "000000000000";
      when "011100000100000" => color_data <= "000000000000";
      when "011100000100001" => color_data <= "000000000000";
      when "011100000100010" => color_data <= "000000000000";
      when "011100000100011" => color_data <= "000000000000";
      when "011100000100100" => color_data <= "000000000000";
      when "011100000100101" => color_data <= "000000000000";
      when "011100000100110" => color_data <= "000000000000";
      when "011100000100111" => color_data <= "000000000000";
      when "011100000101000" => color_data <= "000000000000";
      when "011100000101001" => color_data <= "000000000000";
      when "011100000101010" => color_data <= "000000000000";
      when "011100000101011" => color_data <= "000000000000";
      when "011100000101100" => color_data <= "100001110010";
      when "011100000101101" => color_data <= "111110110000";
      when "011100000101110" => color_data <= "111111000001";
      when "011100000101111" => color_data <= "111111000001";
      when "011100000110000" => color_data <= "111111000001";
      when "011100000110001" => color_data <= "111111000001";
      when "011100000110010" => color_data <= "111111000000";
      when "011100000110011" => color_data <= "111111000000";
      when "011100000110100" => color_data <= "111111000001";
      when "011100000110101" => color_data <= "111111000001";
      when "011100000110110" => color_data <= "111111000001";
      when "011100000110111" => color_data <= "111110110000";
      when "011100000111000" => color_data <= "100101110010";
      when "011100000111001" => color_data <= "000000000000";
      when "011100000111010" => color_data <= "000000000000";
      when "011100000111011" => color_data <= "000000000000";
      when "011100000111100" => color_data <= "000000000000";
      when "011100000111101" => color_data <= "000000000000";
      when "011100000111110" => color_data <= "000000000000";
      when "011100000111111" => color_data <= "000000000000";
      when "011100001000000" => color_data <= "000000000000";
      when "011100001000001" => color_data <= "000000000000";
      when "011100001000010" => color_data <= "000000000000";
      when "011100001000011" => color_data <= "000000000000";
      when "011100001000100" => color_data <= "000000000000";
      when "011100001000101" => color_data <= "000000000000";
      when "011100001000110" => color_data <= "000000000000";
      when "011100001000111" => color_data <= "000000000000";
      when "011100001001000" => color_data <= "000000000000";
      when "011100001001001" => color_data <= "000000000000";
      when "011100001001010" => color_data <= "000000000000";
      when "011100001001011" => color_data <= "000000000000";
      when "011100001001100" => color_data <= "000000000000";
      when "011100001001101" => color_data <= "000000000000";
      when "011100001001110" => color_data <= "000000000000";
      when "011100001001111" => color_data <= "000000000000";
      when "011100001010000" => color_data <= "000000000000";
      when "011100001010001" => color_data <= "000000000000";
      when "011100001010010" => color_data <= "000000000000";
      when "011100001010011" => color_data <= "000000000000";
      when "011100001010100" => color_data <= "000000000000";
      when "011100001010101" => color_data <= "000000000000";
      when "011100001010110" => color_data <= "000000000000";
      when "011100001010111" => color_data <= "000000000000";
      when "011100001011000" => color_data <= "000000000000";
      when "011100001011001" => color_data <= "000000000000";
      when "011100001011010" => color_data <= "000000000000";
      when "011100001011011" => color_data <= "000000000000";
      when "011100001011100" => color_data <= "000000000000";
      when "011100001011101" => color_data <= "000000000000";
      when "011100001011110" => color_data <= "000000000000";
      when "011100001011111" => color_data <= "000000000000";
      when "011100001100000" => color_data <= "000000000000";
      when "011100001100001" => color_data <= "000000000000";
      when "011100001100010" => color_data <= "000000000000";
      when "011100001100011" => color_data <= "000000000000";
      when "011100010000000" => color_data <= "000000000000";
      when "011100010000001" => color_data <= "000000000000";
      when "011100010000010" => color_data <= "000000000000";
      when "011100010000011" => color_data <= "000000000000";
      when "011100010000100" => color_data <= "000000000000";
      when "011100010000101" => color_data <= "000000000000";
      when "011100010000110" => color_data <= "000000000000";
      when "011100010000111" => color_data <= "000000000000";
      when "011100010001000" => color_data <= "000000000000";
      when "011100010001001" => color_data <= "000000000000";
      when "011100010001010" => color_data <= "000000000000";
      when "011100010001011" => color_data <= "000000000000";
      when "011100010001100" => color_data <= "000000000000";
      when "011100010001101" => color_data <= "000000000000";
      when "011100010001110" => color_data <= "000000000000";
      when "011100010001111" => color_data <= "000000000000";
      when "011100010010000" => color_data <= "000000000000";
      when "011100010010001" => color_data <= "000000000000";
      when "011100010010010" => color_data <= "000000000000";
      when "011100010010011" => color_data <= "000000000000";
      when "011100010010100" => color_data <= "000000000000";
      when "011100010010101" => color_data <= "000000000000";
      when "011100010010110" => color_data <= "000000000000";
      when "011100010010111" => color_data <= "000000000000";
      when "011100010011000" => color_data <= "000000000000";
      when "011100010011001" => color_data <= "000000000000";
      when "011100010011010" => color_data <= "000000000000";
      when "011100010011011" => color_data <= "000000000000";
      when "011100010011100" => color_data <= "000000000000";
      when "011100010011101" => color_data <= "000000000000";
      when "011100010011110" => color_data <= "000000000000";
      when "011100010011111" => color_data <= "000000000000";
      when "011100010100000" => color_data <= "000000000000";
      when "011100010100001" => color_data <= "000000000000";
      when "011100010100010" => color_data <= "000000000000";
      when "011100010100011" => color_data <= "000000000000";
      when "011100010100100" => color_data <= "000000000000";
      when "011100010100101" => color_data <= "000000000000";
      when "011100010100110" => color_data <= "000000000000";
      when "011100010100111" => color_data <= "000000000000";
      when "011100010101000" => color_data <= "000000000000";
      when "011100010101001" => color_data <= "000000000000";
      when "011100010101010" => color_data <= "001000100001";
      when "011100010101011" => color_data <= "100110000010";
      when "011100010101100" => color_data <= "110110100000";
      when "011100010101101" => color_data <= "111111000001";
      when "011100010101110" => color_data <= "111111000001";
      when "011100010101111" => color_data <= "111111000001";
      when "011100010110000" => color_data <= "111111000001";
      when "011100010110001" => color_data <= "111111000001";
      when "011100010110010" => color_data <= "111111000001";
      when "011100010110011" => color_data <= "111111000001";
      when "011100010110100" => color_data <= "111111000001";
      when "011100010110101" => color_data <= "111111000001";
      when "011100010110110" => color_data <= "111111000001";
      when "011100010110111" => color_data <= "111111000001";
      when "011100010111000" => color_data <= "110110100000";
      when "011100010111001" => color_data <= "101010000010";
      when "011100010111010" => color_data <= "001100110010";
      when "011100010111011" => color_data <= "000000000000";
      when "011100010111100" => color_data <= "000000000000";
      when "011100010111101" => color_data <= "000000000000";
      when "011100010111110" => color_data <= "000000000000";
      when "011100010111111" => color_data <= "000000000000";
      when "011100011000000" => color_data <= "000000000000";
      when "011100011000001" => color_data <= "000000000000";
      when "011100011000010" => color_data <= "000000000000";
      when "011100011000011" => color_data <= "000000000000";
      when "011100011000100" => color_data <= "000000000000";
      when "011100011000101" => color_data <= "000000000000";
      when "011100011000110" => color_data <= "000000000000";
      when "011100011000111" => color_data <= "000000000000";
      when "011100011001000" => color_data <= "000000000000";
      when "011100011001001" => color_data <= "000000000000";
      when "011100011001010" => color_data <= "000000000000";
      when "011100011001011" => color_data <= "000000000000";
      when "011100011001100" => color_data <= "000000000000";
      when "011100011001101" => color_data <= "000000000000";
      when "011100011001110" => color_data <= "000000000000";
      when "011100011001111" => color_data <= "000000000000";
      when "011100011010000" => color_data <= "000000000000";
      when "011100011010001" => color_data <= "000000000000";
      when "011100011010010" => color_data <= "000000000000";
      when "011100011010011" => color_data <= "000000000000";
      when "011100011010100" => color_data <= "000000000000";
      when "011100011010101" => color_data <= "000000000000";
      when "011100011010110" => color_data <= "000000000000";
      when "011100011010111" => color_data <= "000000000000";
      when "011100011011000" => color_data <= "000000000000";
      when "011100011011001" => color_data <= "000000000000";
      when "011100011011010" => color_data <= "000000000000";
      when "011100011011011" => color_data <= "000000000000";
      when "011100011011100" => color_data <= "000000000000";
      when "011100011011101" => color_data <= "000000000000";
      when "011100011011110" => color_data <= "000000000000";
      when "011100011011111" => color_data <= "000000000000";
      when "011100011100000" => color_data <= "000000000000";
      when "011100011100001" => color_data <= "000000000000";
      when "011100011100010" => color_data <= "000000000000";
      when "011100011100011" => color_data <= "000000000000";
      when "011100100000000" => color_data <= "000000000000";
      when "011100100000001" => color_data <= "000000000000";
      when "011100100000010" => color_data <= "000000000000";
      when "011100100000011" => color_data <= "000000000000";
      when "011100100000100" => color_data <= "000000000000";
      when "011100100000101" => color_data <= "000000000000";
      when "011100100000110" => color_data <= "000000000000";
      when "011100100000111" => color_data <= "000000000000";
      when "011100100001000" => color_data <= "000000000000";
      when "011100100001001" => color_data <= "000000000000";
      when "011100100001010" => color_data <= "000000000000";
      when "011100100001011" => color_data <= "000000000000";
      when "011100100001100" => color_data <= "000000000000";
      when "011100100001101" => color_data <= "000000000000";
      when "011100100001110" => color_data <= "000000000000";
      when "011100100001111" => color_data <= "000000000000";
      when "011100100010000" => color_data <= "000000000000";
      when "011100100010001" => color_data <= "000000000000";
      when "011100100010010" => color_data <= "000000000000";
      when "011100100010011" => color_data <= "000000000000";
      when "011100100010100" => color_data <= "000000000000";
      when "011100100010101" => color_data <= "000000000000";
      when "011100100010110" => color_data <= "000000000000";
      when "011100100010111" => color_data <= "000000000000";
      when "011100100011000" => color_data <= "000000000000";
      when "011100100011001" => color_data <= "000000000000";
      when "011100100011010" => color_data <= "000000000000";
      when "011100100011011" => color_data <= "000000000000";
      when "011100100011100" => color_data <= "000000000000";
      when "011100100011101" => color_data <= "000000000000";
      when "011100100011110" => color_data <= "000000000000";
      when "011100100011111" => color_data <= "000000000000";
      when "011100100100000" => color_data <= "000000000000";
      when "011100100100001" => color_data <= "000000000000";
      when "011100100100010" => color_data <= "000000000000";
      when "011100100100011" => color_data <= "000000000000";
      when "011100100100100" => color_data <= "000000000000";
      when "011100100100101" => color_data <= "000000000000";
      when "011100100100110" => color_data <= "000000000000";
      when "011100100100111" => color_data <= "000000000000";
      when "011100100101000" => color_data <= "000000000000";
      when "011100100101001" => color_data <= "100001110010";
      when "011100100101010" => color_data <= "110110100000";
      when "011100100101011" => color_data <= "111110110000";
      when "011100100101100" => color_data <= "111111000001";
      when "011100100101101" => color_data <= "111111000001";
      when "011100100101110" => color_data <= "111111000001";
      when "011100100101111" => color_data <= "111111000001";
      when "011100100110000" => color_data <= "111111000001";
      when "011100100110001" => color_data <= "111111000001";
      when "011100100110010" => color_data <= "111111000001";
      when "011100100110011" => color_data <= "111111000001";
      when "011100100110100" => color_data <= "111111000001";
      when "011100100110101" => color_data <= "111111000001";
      when "011100100110110" => color_data <= "111111000001";
      when "011100100110111" => color_data <= "111111000001";
      when "011100100111000" => color_data <= "111111000001";
      when "011100100111001" => color_data <= "111110110000";
      when "011100100111010" => color_data <= "110110100000";
      when "011100100111011" => color_data <= "101010000010";
      when "011100100111100" => color_data <= "000100010001";
      when "011100100111101" => color_data <= "000000000000";
      when "011100100111110" => color_data <= "000000000000";
      when "011100100111111" => color_data <= "000000000000";
      when "011100101000000" => color_data <= "000000000000";
      when "011100101000001" => color_data <= "000000000000";
      when "011100101000010" => color_data <= "000000000000";
      when "011100101000011" => color_data <= "000000000000";
      when "011100101000100" => color_data <= "000000000000";
      when "011100101000101" => color_data <= "000000000000";
      when "011100101000110" => color_data <= "000000000000";
      when "011100101000111" => color_data <= "000000000000";
      when "011100101001000" => color_data <= "000000000000";
      when "011100101001001" => color_data <= "000000000000";
      when "011100101001010" => color_data <= "000000000000";
      when "011100101001011" => color_data <= "000000000000";
      when "011100101001100" => color_data <= "000000000000";
      when "011100101001101" => color_data <= "000000000000";
      when "011100101001110" => color_data <= "000000000000";
      when "011100101001111" => color_data <= "000000000000";
      when "011100101010000" => color_data <= "000000000000";
      when "011100101010001" => color_data <= "000000000000";
      when "011100101010010" => color_data <= "000000000000";
      when "011100101010011" => color_data <= "000000000000";
      when "011100101010100" => color_data <= "000000000000";
      when "011100101010101" => color_data <= "000000000000";
      when "011100101010110" => color_data <= "000000000000";
      when "011100101010111" => color_data <= "000000000000";
      when "011100101011000" => color_data <= "000000000000";
      when "011100101011001" => color_data <= "000000000000";
      when "011100101011010" => color_data <= "000000000000";
      when "011100101011011" => color_data <= "000000000000";
      when "011100101011100" => color_data <= "000000000000";
      when "011100101011101" => color_data <= "000000000000";
      when "011100101011110" => color_data <= "000000000000";
      when "011100101011111" => color_data <= "000000000000";
      when "011100101100000" => color_data <= "000000000000";
      when "011100101100001" => color_data <= "000000000000";
      when "011100101100010" => color_data <= "000000000000";
      when "011100101100011" => color_data <= "000000000000";
      when "011100110000000" => color_data <= "000000000000";
      when "011100110000001" => color_data <= "000000000000";
      when "011100110000010" => color_data <= "000000000000";
      when "011100110000011" => color_data <= "000000000000";
      when "011100110000100" => color_data <= "000000000000";
      when "011100110000101" => color_data <= "000000000000";
      when "011100110000110" => color_data <= "000000000000";
      when "011100110000111" => color_data <= "000000000000";
      when "011100110001000" => color_data <= "000000000000";
      when "011100110001001" => color_data <= "000000000000";
      when "011100110001010" => color_data <= "000000000000";
      when "011100110001011" => color_data <= "000000000000";
      when "011100110001100" => color_data <= "000000000000";
      when "011100110001101" => color_data <= "000000000000";
      when "011100110001110" => color_data <= "000000000000";
      when "011100110001111" => color_data <= "000000000000";
      when "011100110010000" => color_data <= "000000000000";
      when "011100110010001" => color_data <= "000000000000";
      when "011100110010010" => color_data <= "000000000000";
      when "011100110010011" => color_data <= "000000000000";
      when "011100110010100" => color_data <= "000000000000";
      when "011100110010101" => color_data <= "000000000000";
      when "011100110010110" => color_data <= "000000000000";
      when "011100110010111" => color_data <= "000000000000";
      when "011100110011000" => color_data <= "000000000000";
      when "011100110011001" => color_data <= "000000000000";
      when "011100110011010" => color_data <= "000000000000";
      when "011100110011011" => color_data <= "000000000000";
      when "011100110011100" => color_data <= "000000000000";
      when "011100110011101" => color_data <= "000000000000";
      when "011100110011110" => color_data <= "000000000000";
      when "011100110011111" => color_data <= "000000000000";
      when "011100110100000" => color_data <= "000000000000";
      when "011100110100001" => color_data <= "000000000000";
      when "011100110100010" => color_data <= "000000000000";
      when "011100110100011" => color_data <= "000000000000";
      when "011100110100100" => color_data <= "000000000000";
      when "011100110100101" => color_data <= "000000000000";
      when "011100110100110" => color_data <= "000000000000";
      when "011100110100111" => color_data <= "001000100001";
      when "011100110101000" => color_data <= "110110100000";
      when "011100110101001" => color_data <= "110110100000";
      when "011100110101010" => color_data <= "111111000000";
      when "011100110101011" => color_data <= "111111000001";
      when "011100110101100" => color_data <= "111111000001";
      when "011100110101101" => color_data <= "111111000001";
      when "011100110101110" => color_data <= "111111000001";
      when "011100110101111" => color_data <= "111111000001";
      when "011100110110000" => color_data <= "111111000001";
      when "011100110110001" => color_data <= "111111000001";
      when "011100110110010" => color_data <= "111111000001";
      when "011100110110011" => color_data <= "111111000001";
      when "011100110110100" => color_data <= "111111000001";
      when "011100110110101" => color_data <= "111111000001";
      when "011100110110110" => color_data <= "111111000001";
      when "011100110110111" => color_data <= "111111000001";
      when "011100110111000" => color_data <= "111111000001";
      when "011100110111001" => color_data <= "111111000001";
      when "011100110111010" => color_data <= "111111000001";
      when "011100110111011" => color_data <= "111110110000";
      when "011100110111100" => color_data <= "110110100000";
      when "011100110111101" => color_data <= "010101000010";
      when "011100110111110" => color_data <= "000000000000";
      when "011100110111111" => color_data <= "000000000000";
      when "011100111000000" => color_data <= "000000000000";
      when "011100111000001" => color_data <= "000000000000";
      when "011100111000010" => color_data <= "000000000000";
      when "011100111000011" => color_data <= "000000000000";
      when "011100111000100" => color_data <= "000000000000";
      when "011100111000101" => color_data <= "000000000000";
      when "011100111000110" => color_data <= "000000000000";
      when "011100111000111" => color_data <= "000000000000";
      when "011100111001000" => color_data <= "000000000000";
      when "011100111001001" => color_data <= "000000000000";
      when "011100111001010" => color_data <= "000000000000";
      when "011100111001011" => color_data <= "000000000000";
      when "011100111001100" => color_data <= "000000000000";
      when "011100111001101" => color_data <= "000000000000";
      when "011100111001110" => color_data <= "000000000000";
      when "011100111001111" => color_data <= "000000000000";
      when "011100111010000" => color_data <= "000000000000";
      when "011100111010001" => color_data <= "000000000000";
      when "011100111010010" => color_data <= "000000000000";
      when "011100111010011" => color_data <= "000000000000";
      when "011100111010100" => color_data <= "000000000000";
      when "011100111010101" => color_data <= "000000000000";
      when "011100111010110" => color_data <= "000000000000";
      when "011100111010111" => color_data <= "000000000000";
      when "011100111011000" => color_data <= "000000000000";
      when "011100111011001" => color_data <= "000000000000";
      when "011100111011010" => color_data <= "000000000000";
      when "011100111011011" => color_data <= "000000000000";
      when "011100111011100" => color_data <= "000000000000";
      when "011100111011101" => color_data <= "000000000000";
      when "011100111011110" => color_data <= "000000000000";
      when "011100111011111" => color_data <= "000000000000";
      when "011100111100000" => color_data <= "000000000000";
      when "011100111100001" => color_data <= "000000000000";
      when "011100111100010" => color_data <= "000000000000";
      when "011100111100011" => color_data <= "000000000000";
      when "011101000000000" => color_data <= "000000000000";
      when "011101000000001" => color_data <= "000000000000";
      when "011101000000010" => color_data <= "000000000000";
      when "011101000000011" => color_data <= "000000000000";
      when "011101000000100" => color_data <= "000000000000";
      when "011101000000101" => color_data <= "000000000000";
      when "011101000000110" => color_data <= "000000000000";
      when "011101000000111" => color_data <= "000000000000";
      when "011101000001000" => color_data <= "000000000000";
      when "011101000001001" => color_data <= "000000000000";
      when "011101000001010" => color_data <= "000000000000";
      when "011101000001011" => color_data <= "000000000000";
      when "011101000001100" => color_data <= "000000000000";
      when "011101000001101" => color_data <= "000000000000";
      when "011101000001110" => color_data <= "000000000000";
      when "011101000001111" => color_data <= "000000000000";
      when "011101000010000" => color_data <= "000000000000";
      when "011101000010001" => color_data <= "000000000000";
      when "011101000010010" => color_data <= "000000000000";
      when "011101000010011" => color_data <= "000000000000";
      when "011101000010100" => color_data <= "000000000000";
      when "011101000010101" => color_data <= "000000000000";
      when "011101000010110" => color_data <= "000000000000";
      when "011101000010111" => color_data <= "000000000000";
      when "011101000011000" => color_data <= "000000000000";
      when "011101000011001" => color_data <= "000000000000";
      when "011101000011010" => color_data <= "000000000000";
      when "011101000011011" => color_data <= "000000000000";
      when "011101000011100" => color_data <= "000000000000";
      when "011101000011101" => color_data <= "000000000000";
      when "011101000011110" => color_data <= "000000000000";
      when "011101000011111" => color_data <= "000000000000";
      when "011101000100000" => color_data <= "000000000000";
      when "011101000100001" => color_data <= "000000000000";
      when "011101000100010" => color_data <= "000000000000";
      when "011101000100011" => color_data <= "000000000000";
      when "011101000100100" => color_data <= "000000000000";
      when "011101000100101" => color_data <= "000000000000";
      when "011101000100110" => color_data <= "000100010001";
      when "011101000100111" => color_data <= "110110100000";
      when "011101000101000" => color_data <= "111110110000";
      when "011101000101001" => color_data <= "111111000001";
      when "011101000101010" => color_data <= "111111000001";
      when "011101000101011" => color_data <= "111111000001";
      when "011101000101100" => color_data <= "111111000001";
      when "011101000101101" => color_data <= "111111000001";
      when "011101000101110" => color_data <= "111111000001";
      when "011101000101111" => color_data <= "111111000001";
      when "011101000110000" => color_data <= "111111000001";
      when "011101000110001" => color_data <= "111111000001";
      when "011101000110010" => color_data <= "111111000001";
      when "011101000110011" => color_data <= "111111000001";
      when "011101000110100" => color_data <= "111111000001";
      when "011101000110101" => color_data <= "111111000001";
      when "011101000110110" => color_data <= "111111000001";
      when "011101000110111" => color_data <= "111111000001";
      when "011101000111000" => color_data <= "111111000001";
      when "011101000111001" => color_data <= "111111000001";
      when "011101000111010" => color_data <= "111111000001";
      when "011101000111011" => color_data <= "111111000001";
      when "011101000111100" => color_data <= "111111000000";
      when "011101000111101" => color_data <= "110110100000";
      when "011101000111110" => color_data <= "010001000010";
      when "011101000111111" => color_data <= "000000000000";
      when "011101001000000" => color_data <= "000000000000";
      when "011101001000001" => color_data <= "000000000000";
      when "011101001000010" => color_data <= "000000000000";
      when "011101001000011" => color_data <= "000000000000";
      when "011101001000100" => color_data <= "000000000000";
      when "011101001000101" => color_data <= "000000000000";
      when "011101001000110" => color_data <= "000000000000";
      when "011101001000111" => color_data <= "000000000000";
      when "011101001001000" => color_data <= "000000000000";
      when "011101001001001" => color_data <= "000000000000";
      when "011101001001010" => color_data <= "000000000000";
      when "011101001001011" => color_data <= "000000000000";
      when "011101001001100" => color_data <= "000000000000";
      when "011101001001101" => color_data <= "000000000000";
      when "011101001001110" => color_data <= "000000000000";
      when "011101001001111" => color_data <= "000000000000";
      when "011101001010000" => color_data <= "000000000000";
      when "011101001010001" => color_data <= "000000000000";
      when "011101001010010" => color_data <= "000000000000";
      when "011101001010011" => color_data <= "000000000000";
      when "011101001010100" => color_data <= "000000000000";
      when "011101001010101" => color_data <= "000000000000";
      when "011101001010110" => color_data <= "000000000000";
      when "011101001010111" => color_data <= "000000000000";
      when "011101001011000" => color_data <= "000000000000";
      when "011101001011001" => color_data <= "000000000000";
      when "011101001011010" => color_data <= "000000000000";
      when "011101001011011" => color_data <= "000000000000";
      when "011101001011100" => color_data <= "000000000000";
      when "011101001011101" => color_data <= "000000000000";
      when "011101001011110" => color_data <= "000000000000";
      when "011101001011111" => color_data <= "000000000000";
      when "011101001100000" => color_data <= "000000000000";
      when "011101001100001" => color_data <= "000000000000";
      when "011101001100010" => color_data <= "000000000000";
      when "011101001100011" => color_data <= "000000000000";
      when "011101010000000" => color_data <= "000000000000";
      when "011101010000001" => color_data <= "000000000000";
      when "011101010000010" => color_data <= "000000000000";
      when "011101010000011" => color_data <= "000000000000";
      when "011101010000100" => color_data <= "000000000000";
      when "011101010000101" => color_data <= "000000000000";
      when "011101010000110" => color_data <= "000000000000";
      when "011101010000111" => color_data <= "000000000000";
      when "011101010001000" => color_data <= "000000000000";
      when "011101010001001" => color_data <= "000000000000";
      when "011101010001010" => color_data <= "000000000000";
      when "011101010001011" => color_data <= "000000000000";
      when "011101010001100" => color_data <= "000000000000";
      when "011101010001101" => color_data <= "000000000000";
      when "011101010001110" => color_data <= "000000000000";
      when "011101010001111" => color_data <= "000000000000";
      when "011101010010000" => color_data <= "000000000000";
      when "011101010010001" => color_data <= "000000000000";
      when "011101010010010" => color_data <= "000000000000";
      when "011101010010011" => color_data <= "000000000000";
      when "011101010010100" => color_data <= "000000000000";
      when "011101010010101" => color_data <= "000000000000";
      when "011101010010110" => color_data <= "000000000000";
      when "011101010010111" => color_data <= "000000000000";
      when "011101010011000" => color_data <= "000000000000";
      when "011101010011001" => color_data <= "000000000000";
      when "011101010011010" => color_data <= "000000000000";
      when "011101010011011" => color_data <= "000000000000";
      when "011101010011100" => color_data <= "000000000000";
      when "011101010011101" => color_data <= "000000000000";
      when "011101010011110" => color_data <= "000000000000";
      when "011101010011111" => color_data <= "000000000000";
      when "011101010100000" => color_data <= "000000000000";
      when "011101010100001" => color_data <= "000000000000";
      when "011101010100010" => color_data <= "000000000000";
      when "011101010100011" => color_data <= "000000000000";
      when "011101010100100" => color_data <= "000000000000";
      when "011101010100101" => color_data <= "000000000000";
      when "011101010100110" => color_data <= "110010100000";
      when "011101010100111" => color_data <= "111110110000";
      when "011101010101000" => color_data <= "111111000001";
      when "011101010101001" => color_data <= "111111000001";
      when "011101010101010" => color_data <= "111111000001";
      when "011101010101011" => color_data <= "111111000001";
      when "011101010101100" => color_data <= "111111000001";
      when "011101010101101" => color_data <= "111111000001";
      when "011101010101110" => color_data <= "111111000001";
      when "011101010101111" => color_data <= "111111000001";
      when "011101010110000" => color_data <= "111111000001";
      when "011101010110001" => color_data <= "111111000001";
      when "011101010110010" => color_data <= "111111000001";
      when "011101010110011" => color_data <= "111111000001";
      when "011101010110100" => color_data <= "111111000001";
      when "011101010110101" => color_data <= "111111000001";
      when "011101010110110" => color_data <= "111111000001";
      when "011101010110111" => color_data <= "111111000001";
      when "011101010111000" => color_data <= "111111000001";
      when "011101010111001" => color_data <= "111111000001";
      when "011101010111010" => color_data <= "111111000001";
      when "011101010111011" => color_data <= "111111000001";
      when "011101010111100" => color_data <= "111111000001";
      when "011101010111101" => color_data <= "111111000000";
      when "011101010111110" => color_data <= "110110100000";
      when "011101010111111" => color_data <= "000100010001";
      when "011101011000000" => color_data <= "000000000000";
      when "011101011000001" => color_data <= "000000000000";
      when "011101011000010" => color_data <= "000000000000";
      when "011101011000011" => color_data <= "000000000000";
      when "011101011000100" => color_data <= "000000000000";
      when "011101011000101" => color_data <= "000000000000";
      when "011101011000110" => color_data <= "000000000000";
      when "011101011000111" => color_data <= "000000000000";
      when "011101011001000" => color_data <= "000000000000";
      when "011101011001001" => color_data <= "000000000000";
      when "011101011001010" => color_data <= "000000000000";
      when "011101011001011" => color_data <= "000000000000";
      when "011101011001100" => color_data <= "000000000000";
      when "011101011001101" => color_data <= "000000000000";
      when "011101011001110" => color_data <= "000000000000";
      when "011101011001111" => color_data <= "000000000000";
      when "011101011010000" => color_data <= "000000000000";
      when "011101011010001" => color_data <= "000000000000";
      when "011101011010010" => color_data <= "000000000000";
      when "011101011010011" => color_data <= "000000000000";
      when "011101011010100" => color_data <= "000000000000";
      when "011101011010101" => color_data <= "000000000000";
      when "011101011010110" => color_data <= "000000000000";
      when "011101011010111" => color_data <= "000000000000";
      when "011101011011000" => color_data <= "000000000000";
      when "011101011011001" => color_data <= "000000000000";
      when "011101011011010" => color_data <= "000000000000";
      when "011101011011011" => color_data <= "000000000000";
      when "011101011011100" => color_data <= "000000000000";
      when "011101011011101" => color_data <= "000000000000";
      when "011101011011110" => color_data <= "000000000000";
      when "011101011011111" => color_data <= "000000000000";
      when "011101011100000" => color_data <= "000000000000";
      when "011101011100001" => color_data <= "000000000000";
      when "011101011100010" => color_data <= "000000000000";
      when "011101011100011" => color_data <= "000000000000";
      when "011101100000000" => color_data <= "000000000000";
      when "011101100000001" => color_data <= "000000000000";
      when "011101100000010" => color_data <= "000000000000";
      when "011101100000011" => color_data <= "000000000000";
      when "011101100000100" => color_data <= "000000000000";
      when "011101100000101" => color_data <= "000000000000";
      when "011101100000110" => color_data <= "000000000000";
      when "011101100000111" => color_data <= "000000000000";
      when "011101100001000" => color_data <= "000000000000";
      when "011101100001001" => color_data <= "000000000000";
      when "011101100001010" => color_data <= "000000000000";
      when "011101100001011" => color_data <= "000000000000";
      when "011101100001100" => color_data <= "000000000000";
      when "011101100001101" => color_data <= "000000000000";
      when "011101100001110" => color_data <= "000000000000";
      when "011101100001111" => color_data <= "000000000000";
      when "011101100010000" => color_data <= "000000000000";
      when "011101100010001" => color_data <= "000000000000";
      when "011101100010010" => color_data <= "000000000000";
      when "011101100010011" => color_data <= "000000000000";
      when "011101100010100" => color_data <= "000000000000";
      when "011101100010101" => color_data <= "000000000000";
      when "011101100010110" => color_data <= "000000000000";
      when "011101100010111" => color_data <= "000000000000";
      when "011101100011000" => color_data <= "000000000000";
      when "011101100011001" => color_data <= "000000000000";
      when "011101100011010" => color_data <= "000000000000";
      when "011101100011011" => color_data <= "000000000000";
      when "011101100011100" => color_data <= "000000000000";
      when "011101100011101" => color_data <= "000000000000";
      when "011101100011110" => color_data <= "000000000000";
      when "011101100011111" => color_data <= "000000000000";
      when "011101100100000" => color_data <= "000000000000";
      when "011101100100001" => color_data <= "000000000000";
      when "011101100100010" => color_data <= "000000000000";
      when "011101100100011" => color_data <= "000000000000";
      when "011101100100100" => color_data <= "000000000000";
      when "011101100100101" => color_data <= "011001010011";
      when "011101100100110" => color_data <= "110110100000";
      when "011101100100111" => color_data <= "111111000001";
      when "011101100101000" => color_data <= "111111000001";
      when "011101100101001" => color_data <= "111111000001";
      when "011101100101010" => color_data <= "111111000001";
      when "011101100101011" => color_data <= "111111000001";
      when "011101100101100" => color_data <= "111111000001";
      when "011101100101101" => color_data <= "111111000001";
      when "011101100101110" => color_data <= "111111000001";
      when "011101100101111" => color_data <= "111111000001";
      when "011101100110000" => color_data <= "111111000001";
      when "011101100110001" => color_data <= "111111000001";
      when "011101100110010" => color_data <= "111111000001";
      when "011101100110011" => color_data <= "111111000001";
      when "011101100110100" => color_data <= "111111000001";
      when "011101100110101" => color_data <= "111111000001";
      when "011101100110110" => color_data <= "111111000001";
      when "011101100110111" => color_data <= "111111000001";
      when "011101100111000" => color_data <= "111111000001";
      when "011101100111001" => color_data <= "111111000001";
      when "011101100111010" => color_data <= "111111000001";
      when "011101100111011" => color_data <= "111111000001";
      when "011101100111100" => color_data <= "111111000001";
      when "011101100111101" => color_data <= "111111000001";
      when "011101100111110" => color_data <= "111110110000";
      when "011101100111111" => color_data <= "100110000010";
      when "011101101000000" => color_data <= "000000000000";
      when "011101101000001" => color_data <= "000000000000";
      when "011101101000010" => color_data <= "000000000000";
      when "011101101000011" => color_data <= "000000000000";
      when "011101101000100" => color_data <= "000000000000";
      when "011101101000101" => color_data <= "000000000000";
      when "011101101000110" => color_data <= "000000000000";
      when "011101101000111" => color_data <= "000000000000";
      when "011101101001000" => color_data <= "000000000000";
      when "011101101001001" => color_data <= "000000000000";
      when "011101101001010" => color_data <= "000000000000";
      when "011101101001011" => color_data <= "000000000000";
      when "011101101001100" => color_data <= "000000000000";
      when "011101101001101" => color_data <= "000000000000";
      when "011101101001110" => color_data <= "000000000000";
      when "011101101001111" => color_data <= "000000000000";
      when "011101101010000" => color_data <= "000000000000";
      when "011101101010001" => color_data <= "000000000000";
      when "011101101010010" => color_data <= "000000000000";
      when "011101101010011" => color_data <= "000000000000";
      when "011101101010100" => color_data <= "000000000000";
      when "011101101010101" => color_data <= "000000000000";
      when "011101101010110" => color_data <= "000000000000";
      when "011101101010111" => color_data <= "000000000000";
      when "011101101011000" => color_data <= "000000000000";
      when "011101101011001" => color_data <= "000000000000";
      when "011101101011010" => color_data <= "000000000000";
      when "011101101011011" => color_data <= "000000000000";
      when "011101101011100" => color_data <= "000000000000";
      when "011101101011101" => color_data <= "000000000000";
      when "011101101011110" => color_data <= "000000000000";
      when "011101101011111" => color_data <= "000000000000";
      when "011101101100000" => color_data <= "000000000000";
      when "011101101100001" => color_data <= "000000000000";
      when "011101101100010" => color_data <= "000000000000";
      when "011101101100011" => color_data <= "000000000000";
      when "011101110000000" => color_data <= "000000000000";
      when "011101110000001" => color_data <= "000000000000";
      when "011101110000010" => color_data <= "000000000000";
      when "011101110000011" => color_data <= "000000000000";
      when "011101110000100" => color_data <= "000000000000";
      when "011101110000101" => color_data <= "000000000000";
      when "011101110000110" => color_data <= "000000000000";
      when "011101110000111" => color_data <= "000000000000";
      when "011101110001000" => color_data <= "000000000000";
      when "011101110001001" => color_data <= "000000000000";
      when "011101110001010" => color_data <= "000000000000";
      when "011101110001011" => color_data <= "000000000000";
      when "011101110001100" => color_data <= "000000000000";
      when "011101110001101" => color_data <= "000000000000";
      when "011101110001110" => color_data <= "000000000000";
      when "011101110001111" => color_data <= "000000000000";
      when "011101110010000" => color_data <= "000000000000";
      when "011101110010001" => color_data <= "000000000000";
      when "011101110010010" => color_data <= "000000000000";
      when "011101110010011" => color_data <= "000000000000";
      when "011101110010100" => color_data <= "000000000000";
      when "011101110010101" => color_data <= "000000000000";
      when "011101110010110" => color_data <= "000000000000";
      when "011101110010111" => color_data <= "000000000000";
      when "011101110011000" => color_data <= "000000000000";
      when "011101110011001" => color_data <= "000000000000";
      when "011101110011010" => color_data <= "000000000000";
      when "011101110011011" => color_data <= "000000000000";
      when "011101110011100" => color_data <= "000000000000";
      when "011101110011101" => color_data <= "000000000000";
      when "011101110011110" => color_data <= "000000000000";
      when "011101110011111" => color_data <= "000000000000";
      when "011101110100000" => color_data <= "000000000000";
      when "011101110100001" => color_data <= "000000000000";
      when "011101110100010" => color_data <= "000000000000";
      when "011101110100011" => color_data <= "000000000000";
      when "011101110100100" => color_data <= "000000000000";
      when "011101110100101" => color_data <= "110010010001";
      when "011101110100110" => color_data <= "111111000000";
      when "011101110100111" => color_data <= "111111000001";
      when "011101110101000" => color_data <= "111111000001";
      when "011101110101001" => color_data <= "111111000001";
      when "011101110101010" => color_data <= "111111000001";
      when "011101110101011" => color_data <= "111111000001";
      when "011101110101100" => color_data <= "111111000001";
      when "011101110101101" => color_data <= "111111000001";
      when "011101110101110" => color_data <= "111111000001";
      when "011101110101111" => color_data <= "111111000001";
      when "011101110110000" => color_data <= "111111000001";
      when "011101110110001" => color_data <= "111111000001";
      when "011101110110010" => color_data <= "111111000001";
      when "011101110110011" => color_data <= "111111000001";
      when "011101110110100" => color_data <= "111111000001";
      when "011101110110101" => color_data <= "111111000001";
      when "011101110110110" => color_data <= "111111000001";
      when "011101110110111" => color_data <= "111111000001";
      when "011101110111000" => color_data <= "111111000001";
      when "011101110111001" => color_data <= "111111000001";
      when "011101110111010" => color_data <= "111111000001";
      when "011101110111011" => color_data <= "111111000001";
      when "011101110111100" => color_data <= "111111000001";
      when "011101110111101" => color_data <= "111111000001";
      when "011101110111110" => color_data <= "111111000000";
      when "011101110111111" => color_data <= "110110100000";
      when "011101111000000" => color_data <= "000100010001";
      when "011101111000001" => color_data <= "000000000000";
      when "011101111000010" => color_data <= "000000000000";
      when "011101111000011" => color_data <= "000000000000";
      when "011101111000100" => color_data <= "000000000000";
      when "011101111000101" => color_data <= "000000000000";
      when "011101111000110" => color_data <= "000000000000";
      when "011101111000111" => color_data <= "000000000000";
      when "011101111001000" => color_data <= "000000000000";
      when "011101111001001" => color_data <= "000000000000";
      when "011101111001010" => color_data <= "000000000000";
      when "011101111001011" => color_data <= "000000000000";
      when "011101111001100" => color_data <= "000000000000";
      when "011101111001101" => color_data <= "000000000000";
      when "011101111001110" => color_data <= "000000000000";
      when "011101111001111" => color_data <= "000000000000";
      when "011101111010000" => color_data <= "000000000000";
      when "011101111010001" => color_data <= "000000000000";
      when "011101111010010" => color_data <= "000000000000";
      when "011101111010011" => color_data <= "000000000000";
      when "011101111010100" => color_data <= "000000000000";
      when "011101111010101" => color_data <= "000000000000";
      when "011101111010110" => color_data <= "000000000000";
      when "011101111010111" => color_data <= "000000000000";
      when "011101111011000" => color_data <= "000000000000";
      when "011101111011001" => color_data <= "000000000000";
      when "011101111011010" => color_data <= "000000000000";
      when "011101111011011" => color_data <= "000000000000";
      when "011101111011100" => color_data <= "000000000000";
      when "011101111011101" => color_data <= "000000000000";
      when "011101111011110" => color_data <= "000000000000";
      when "011101111011111" => color_data <= "000000000000";
      when "011101111100000" => color_data <= "000000000000";
      when "011101111100001" => color_data <= "000000000000";
      when "011101111100010" => color_data <= "000000000000";
      when "011101111100011" => color_data <= "000000000000";
      when "011110000000000" => color_data <= "000000000000";
      when "011110000000001" => color_data <= "000000000000";
      when "011110000000010" => color_data <= "000000000000";
      when "011110000000011" => color_data <= "000000000000";
      when "011110000000100" => color_data <= "000000000000";
      when "011110000000101" => color_data <= "000000000000";
      when "011110000000110" => color_data <= "000000000000";
      when "011110000000111" => color_data <= "000000000000";
      when "011110000001000" => color_data <= "000000000000";
      when "011110000001001" => color_data <= "000000000000";
      when "011110000001010" => color_data <= "000000000000";
      when "011110000001011" => color_data <= "000000000000";
      when "011110000001100" => color_data <= "000000000000";
      when "011110000001101" => color_data <= "000000000000";
      when "011110000001110" => color_data <= "000000000000";
      when "011110000001111" => color_data <= "000000000000";
      when "011110000010000" => color_data <= "000000000000";
      when "011110000010001" => color_data <= "000000000000";
      when "011110000010010" => color_data <= "000000000000";
      when "011110000010011" => color_data <= "000000000000";
      when "011110000010100" => color_data <= "000000000000";
      when "011110000010101" => color_data <= "000000000000";
      when "011110000010110" => color_data <= "000000000000";
      when "011110000010111" => color_data <= "000000000000";
      when "011110000011000" => color_data <= "000000000000";
      when "011110000011001" => color_data <= "000000000000";
      when "011110000011010" => color_data <= "000000000000";
      when "011110000011011" => color_data <= "000000000000";
      when "011110000011100" => color_data <= "000000000000";
      when "011110000011101" => color_data <= "000000000000";
      when "011110000011110" => color_data <= "000000000000";
      when "011110000011111" => color_data <= "000000000000";
      when "011110000100000" => color_data <= "000000000000";
      when "011110000100001" => color_data <= "000000000000";
      when "011110000100010" => color_data <= "000000000000";
      when "011110000100011" => color_data <= "000000000000";
      when "011110000100100" => color_data <= "001100100010";
      when "011110000100101" => color_data <= "110110100000";
      when "011110000100110" => color_data <= "111111000001";
      when "011110000100111" => color_data <= "111111000001";
      when "011110000101000" => color_data <= "111111000001";
      when "011110000101001" => color_data <= "111111000001";
      when "011110000101010" => color_data <= "111111000001";
      when "011110000101011" => color_data <= "111111000001";
      when "011110000101100" => color_data <= "111111000001";
      when "011110000101101" => color_data <= "111111000001";
      when "011110000101110" => color_data <= "111111000001";
      when "011110000101111" => color_data <= "111111000001";
      when "011110000110000" => color_data <= "111111000001";
      when "011110000110001" => color_data <= "111111000001";
      when "011110000110010" => color_data <= "111111000001";
      when "011110000110011" => color_data <= "111111000001";
      when "011110000110100" => color_data <= "111111000001";
      when "011110000110101" => color_data <= "111111000001";
      when "011110000110110" => color_data <= "111111000001";
      when "011110000110111" => color_data <= "111111000001";
      when "011110000111000" => color_data <= "111111000001";
      when "011110000111001" => color_data <= "111111000001";
      when "011110000111010" => color_data <= "111111000001";
      when "011110000111011" => color_data <= "111111000001";
      when "011110000111100" => color_data <= "111111000001";
      when "011110000111101" => color_data <= "111111000001";
      when "011110000111110" => color_data <= "111111000001";
      when "011110000111111" => color_data <= "111110110000";
      when "011110001000000" => color_data <= "010101010011";
      when "011110001000001" => color_data <= "000000000000";
      when "011110001000010" => color_data <= "000000000000";
      when "011110001000011" => color_data <= "000000000000";
      when "011110001000100" => color_data <= "000000000000";
      when "011110001000101" => color_data <= "000000000000";
      when "011110001000110" => color_data <= "000000000000";
      when "011110001000111" => color_data <= "000000000000";
      when "011110001001000" => color_data <= "000000000000";
      when "011110001001001" => color_data <= "000000000000";
      when "011110001001010" => color_data <= "000000000000";
      when "011110001001011" => color_data <= "000000000000";
      when "011110001001100" => color_data <= "000000000000";
      when "011110001001101" => color_data <= "000000000000";
      when "011110001001110" => color_data <= "000000000000";
      when "011110001001111" => color_data <= "000000000000";
      when "011110001010000" => color_data <= "000000000000";
      when "011110001010001" => color_data <= "000000000000";
      when "011110001010010" => color_data <= "000000000000";
      when "011110001010011" => color_data <= "000000000000";
      when "011110001010100" => color_data <= "000000000000";
      when "011110001010101" => color_data <= "000000000000";
      when "011110001010110" => color_data <= "000000000000";
      when "011110001010111" => color_data <= "000000000000";
      when "011110001011000" => color_data <= "000000000000";
      when "011110001011001" => color_data <= "000000000000";
      when "011110001011010" => color_data <= "000000000000";
      when "011110001011011" => color_data <= "000000000000";
      when "011110001011100" => color_data <= "000000000000";
      when "011110001011101" => color_data <= "000000000000";
      when "011110001011110" => color_data <= "000000000000";
      when "011110001011111" => color_data <= "000000000000";
      when "011110001100000" => color_data <= "000000000000";
      when "011110001100001" => color_data <= "000000000000";
      when "011110001100010" => color_data <= "000000000000";
      when "011110001100011" => color_data <= "000000000000";
      when "011110010000000" => color_data <= "000000000000";
      when "011110010000001" => color_data <= "000000000000";
      when "011110010000010" => color_data <= "000000000000";
      when "011110010000011" => color_data <= "000000000000";
      when "011110010000100" => color_data <= "000000000000";
      when "011110010000101" => color_data <= "000000000000";
      when "011110010000110" => color_data <= "000000000000";
      when "011110010000111" => color_data <= "000000000000";
      when "011110010001000" => color_data <= "000000000000";
      when "011110010001001" => color_data <= "000000000000";
      when "011110010001010" => color_data <= "000000000000";
      when "011110010001011" => color_data <= "000000000000";
      when "011110010001100" => color_data <= "000000000000";
      when "011110010001101" => color_data <= "000000000000";
      when "011110010001110" => color_data <= "000000000000";
      when "011110010001111" => color_data <= "000000000000";
      when "011110010010000" => color_data <= "000000000000";
      when "011110010010001" => color_data <= "000000000000";
      when "011110010010010" => color_data <= "000000000000";
      when "011110010010011" => color_data <= "000000000000";
      when "011110010010100" => color_data <= "000000000000";
      when "011110010010101" => color_data <= "000000000000";
      when "011110010010110" => color_data <= "000000000000";
      when "011110010010111" => color_data <= "000000000000";
      when "011110010011000" => color_data <= "000000000000";
      when "011110010011001" => color_data <= "000000000000";
      when "011110010011010" => color_data <= "000000000000";
      when "011110010011011" => color_data <= "000000000000";
      when "011110010011100" => color_data <= "000000000000";
      when "011110010011101" => color_data <= "000000000000";
      when "011110010011110" => color_data <= "000000000000";
      when "011110010011111" => color_data <= "000000000000";
      when "011110010100000" => color_data <= "000000000000";
      when "011110010100001" => color_data <= "000000000000";
      when "011110010100010" => color_data <= "000000000000";
      when "011110010100011" => color_data <= "000000000000";
      when "011110010100100" => color_data <= "001100110010";
      when "011110010100101" => color_data <= "111110110000";
      when "011110010100110" => color_data <= "111111000001";
      when "011110010100111" => color_data <= "111111000001";
      when "011110010101000" => color_data <= "111111000001";
      when "011110010101001" => color_data <= "111111000001";
      when "011110010101010" => color_data <= "111111000001";
      when "011110010101011" => color_data <= "111111000001";
      when "011110010101100" => color_data <= "111111000001";
      when "011110010101101" => color_data <= "111111000001";
      when "011110010101110" => color_data <= "111111000001";
      when "011110010101111" => color_data <= "111111000001";
      when "011110010110000" => color_data <= "111111000001";
      when "011110010110001" => color_data <= "111111000001";
      when "011110010110010" => color_data <= "111111000001";
      when "011110010110011" => color_data <= "111111000001";
      when "011110010110100" => color_data <= "111111000001";
      when "011110010110101" => color_data <= "111111000001";
      when "011110010110110" => color_data <= "111111000001";
      when "011110010110111" => color_data <= "111111000001";
      when "011110010111000" => color_data <= "111111000001";
      when "011110010111001" => color_data <= "111111000001";
      when "011110010111010" => color_data <= "111111000001";
      when "011110010111011" => color_data <= "111111000001";
      when "011110010111100" => color_data <= "111111000001";
      when "011110010111101" => color_data <= "111111000001";
      when "011110010111110" => color_data <= "111111000001";
      when "011110010111111" => color_data <= "111110110000";
      when "011110011000000" => color_data <= "011001100011";
      when "011110011000001" => color_data <= "000000000000";
      when "011110011000010" => color_data <= "000000000000";
      when "011110011000011" => color_data <= "000000000000";
      when "011110011000100" => color_data <= "000000000000";
      when "011110011000101" => color_data <= "000000000000";
      when "011110011000110" => color_data <= "000000000000";
      when "011110011000111" => color_data <= "000000000000";
      when "011110011001000" => color_data <= "000000000000";
      when "011110011001001" => color_data <= "000000000000";
      when "011110011001010" => color_data <= "000000000000";
      when "011110011001011" => color_data <= "000000000000";
      when "011110011001100" => color_data <= "000000000000";
      when "011110011001101" => color_data <= "000000000000";
      when "011110011001110" => color_data <= "000000000000";
      when "011110011001111" => color_data <= "000000000000";
      when "011110011010000" => color_data <= "000000000000";
      when "011110011010001" => color_data <= "000000000000";
      when "011110011010010" => color_data <= "000000000000";
      when "011110011010011" => color_data <= "000000000000";
      when "011110011010100" => color_data <= "000000000000";
      when "011110011010101" => color_data <= "000000000000";
      when "011110011010110" => color_data <= "000000000000";
      when "011110011010111" => color_data <= "000000000000";
      when "011110011011000" => color_data <= "000000000000";
      when "011110011011001" => color_data <= "000000000000";
      when "011110011011010" => color_data <= "000000000000";
      when "011110011011011" => color_data <= "000000000000";
      when "011110011011100" => color_data <= "000000000000";
      when "011110011011101" => color_data <= "000000000000";
      when "011110011011110" => color_data <= "000000000000";
      when "011110011011111" => color_data <= "000000000000";
      when "011110011100000" => color_data <= "000000000000";
      when "011110011100001" => color_data <= "000000000000";
      when "011110011100010" => color_data <= "000000000000";
      when "011110011100011" => color_data <= "000000000000";
      when "011110100000000" => color_data <= "000000000000";
      when "011110100000001" => color_data <= "000000000000";
      when "011110100000010" => color_data <= "000000000000";
      when "011110100000011" => color_data <= "000000000000";
      when "011110100000100" => color_data <= "000000000000";
      when "011110100000101" => color_data <= "000000000000";
      when "011110100000110" => color_data <= "000000000000";
      when "011110100000111" => color_data <= "000000000000";
      when "011110100001000" => color_data <= "000000000000";
      when "011110100001001" => color_data <= "000000000000";
      when "011110100001010" => color_data <= "000000000000";
      when "011110100001011" => color_data <= "000000000000";
      when "011110100001100" => color_data <= "000000000000";
      when "011110100001101" => color_data <= "000000000000";
      when "011110100001110" => color_data <= "000000000000";
      when "011110100001111" => color_data <= "000000000000";
      when "011110100010000" => color_data <= "000000000000";
      when "011110100010001" => color_data <= "000000000000";
      when "011110100010010" => color_data <= "000000000000";
      when "011110100010011" => color_data <= "000000000000";
      when "011110100010100" => color_data <= "000000000000";
      when "011110100010101" => color_data <= "000000000000";
      when "011110100010110" => color_data <= "000000000000";
      when "011110100010111" => color_data <= "000000000000";
      when "011110100011000" => color_data <= "000000000000";
      when "011110100011001" => color_data <= "000000000000";
      when "011110100011010" => color_data <= "000000000000";
      when "011110100011011" => color_data <= "000000000000";
      when "011110100011100" => color_data <= "000000000000";
      when "011110100011101" => color_data <= "000000000000";
      when "011110100011110" => color_data <= "000000000000";
      when "011110100011111" => color_data <= "000000000000";
      when "011110100100000" => color_data <= "000000000000";
      when "011110100100001" => color_data <= "000000000000";
      when "011110100100010" => color_data <= "000100010001";
      when "011110100100011" => color_data <= "000000000000";
      when "011110100100100" => color_data <= "011001010011";
      when "011110100100101" => color_data <= "111110110000";
      when "011110100100110" => color_data <= "111111000001";
      when "011110100100111" => color_data <= "111111000001";
      when "011110100101000" => color_data <= "111111000001";
      when "011110100101001" => color_data <= "111111000001";
      when "011110100101010" => color_data <= "111111000001";
      when "011110100101011" => color_data <= "111111000001";
      when "011110100101100" => color_data <= "111111000001";
      when "011110100101101" => color_data <= "111111000001";
      when "011110100101110" => color_data <= "111111000001";
      when "011110100101111" => color_data <= "111111000001";
      when "011110100110000" => color_data <= "111111000001";
      when "011110100110001" => color_data <= "111111000001";
      when "011110100110010" => color_data <= "111111000001";
      when "011110100110011" => color_data <= "111111000001";
      when "011110100110100" => color_data <= "111111000001";
      when "011110100110101" => color_data <= "111111000001";
      when "011110100110110" => color_data <= "111111000001";
      when "011110100110111" => color_data <= "111111000001";
      when "011110100111000" => color_data <= "111111000001";
      when "011110100111001" => color_data <= "111111000001";
      when "011110100111010" => color_data <= "111111000001";
      when "011110100111011" => color_data <= "111111000001";
      when "011110100111100" => color_data <= "111111000001";
      when "011110100111101" => color_data <= "111111000001";
      when "011110100111110" => color_data <= "111111000001";
      when "011110100111111" => color_data <= "111110110000";
      when "011110101000000" => color_data <= "100001110010";
      when "011110101000001" => color_data <= "000000000000";
      when "011110101000010" => color_data <= "000100010000";
      when "011110101000011" => color_data <= "000000000000";
      when "011110101000100" => color_data <= "000000000000";
      when "011110101000101" => color_data <= "000000000000";
      when "011110101000110" => color_data <= "000000000000";
      when "011110101000111" => color_data <= "000000000000";
      when "011110101001000" => color_data <= "000000000000";
      when "011110101001001" => color_data <= "000000000000";
      when "011110101001010" => color_data <= "000000000000";
      when "011110101001011" => color_data <= "000000000000";
      when "011110101001100" => color_data <= "000000000000";
      when "011110101001101" => color_data <= "000000000000";
      when "011110101001110" => color_data <= "000000000000";
      when "011110101001111" => color_data <= "000000000000";
      when "011110101010000" => color_data <= "000000000000";
      when "011110101010001" => color_data <= "000000000000";
      when "011110101010010" => color_data <= "000000000000";
      when "011110101010011" => color_data <= "000000000000";
      when "011110101010100" => color_data <= "000000000000";
      when "011110101010101" => color_data <= "000000000000";
      when "011110101010110" => color_data <= "000000000000";
      when "011110101010111" => color_data <= "000000000000";
      when "011110101011000" => color_data <= "000000000000";
      when "011110101011001" => color_data <= "000000000000";
      when "011110101011010" => color_data <= "000000000000";
      when "011110101011011" => color_data <= "000000000000";
      when "011110101011100" => color_data <= "000000000000";
      when "011110101011101" => color_data <= "000000000000";
      when "011110101011110" => color_data <= "000000000000";
      when "011110101011111" => color_data <= "000000000000";
      when "011110101100000" => color_data <= "000000000000";
      when "011110101100001" => color_data <= "000000000000";
      when "011110101100010" => color_data <= "000000000000";
      when "011110101100011" => color_data <= "000000000000";
      when "011110110000000" => color_data <= "000000000000";
      when "011110110000001" => color_data <= "000000000000";
      when "011110110000010" => color_data <= "000000000000";
      when "011110110000011" => color_data <= "000000000000";
      when "011110110000100" => color_data <= "000000000000";
      when "011110110000101" => color_data <= "000000000000";
      when "011110110000110" => color_data <= "000000000000";
      when "011110110000111" => color_data <= "000000000000";
      when "011110110001000" => color_data <= "000000000000";
      when "011110110001001" => color_data <= "000000000000";
      when "011110110001010" => color_data <= "000000000000";
      when "011110110001011" => color_data <= "000000000000";
      when "011110110001100" => color_data <= "000000000000";
      when "011110110001101" => color_data <= "000000000000";
      when "011110110001110" => color_data <= "000000000000";
      when "011110110001111" => color_data <= "000000000000";
      when "011110110010000" => color_data <= "000000000000";
      when "011110110010001" => color_data <= "000000000000";
      when "011110110010010" => color_data <= "000000000000";
      when "011110110010011" => color_data <= "000000000000";
      when "011110110010100" => color_data <= "000000000000";
      when "011110110010101" => color_data <= "000000000000";
      when "011110110010110" => color_data <= "000000000000";
      when "011110110010111" => color_data <= "000000000000";
      when "011110110011000" => color_data <= "000000000000";
      when "011110110011001" => color_data <= "000000000000";
      when "011110110011010" => color_data <= "000000000000";
      when "011110110011011" => color_data <= "000000000000";
      when "011110110011100" => color_data <= "000000000000";
      when "011110110011101" => color_data <= "000000000000";
      when "011110110011110" => color_data <= "000000000000";
      when "011110110011111" => color_data <= "000000000000";
      when "011110110100000" => color_data <= "000000000000";
      when "011110110100001" => color_data <= "010101010011";
      when "011110110100010" => color_data <= "110110100000";
      when "011110110100011" => color_data <= "111111000000";
      when "011110110100100" => color_data <= "111111000001";
      when "011110110100101" => color_data <= "111111000001";
      when "011110110100110" => color_data <= "111111000001";
      when "011110110100111" => color_data <= "111111000001";
      when "011110110101000" => color_data <= "111111000001";
      when "011110110101001" => color_data <= "111111000001";
      when "011110110101010" => color_data <= "111111000001";
      when "011110110101011" => color_data <= "111111000001";
      when "011110110101100" => color_data <= "111111000001";
      when "011110110101101" => color_data <= "111111000001";
      when "011110110101110" => color_data <= "111111000001";
      when "011110110101111" => color_data <= "111111000001";
      when "011110110110000" => color_data <= "111111000001";
      when "011110110110001" => color_data <= "111111000001";
      when "011110110110010" => color_data <= "111111000001";
      when "011110110110011" => color_data <= "111111000001";
      when "011110110110100" => color_data <= "111111000001";
      when "011110110110101" => color_data <= "111111000001";
      when "011110110110110" => color_data <= "111111000001";
      when "011110110110111" => color_data <= "111111000001";
      when "011110110111000" => color_data <= "111111000001";
      when "011110110111001" => color_data <= "111111000001";
      when "011110110111010" => color_data <= "111111000001";
      when "011110110111011" => color_data <= "111111000001";
      when "011110110111100" => color_data <= "111111000001";
      when "011110110111101" => color_data <= "111111000001";
      when "011110110111110" => color_data <= "111111000001";
      when "011110110111111" => color_data <= "111111000001";
      when "011110111000000" => color_data <= "111111000000";
      when "011110111000001" => color_data <= "111111000000";
      when "011110111000010" => color_data <= "111110110000";
      when "011110111000011" => color_data <= "100001110010";
      when "011110111000100" => color_data <= "000000000000";
      when "011110111000101" => color_data <= "000000000000";
      when "011110111000110" => color_data <= "000000000000";
      when "011110111000111" => color_data <= "000000000000";
      when "011110111001000" => color_data <= "000000000000";
      when "011110111001001" => color_data <= "000000000000";
      when "011110111001010" => color_data <= "000000000000";
      when "011110111001011" => color_data <= "000000000000";
      when "011110111001100" => color_data <= "000000000000";
      when "011110111001101" => color_data <= "000000000000";
      when "011110111001110" => color_data <= "000000000000";
      when "011110111001111" => color_data <= "000000000000";
      when "011110111010000" => color_data <= "000000000000";
      when "011110111010001" => color_data <= "000000000000";
      when "011110111010010" => color_data <= "000000000000";
      when "011110111010011" => color_data <= "000000000000";
      when "011110111010100" => color_data <= "000000000000";
      when "011110111010101" => color_data <= "000000000000";
      when "011110111010110" => color_data <= "000000000000";
      when "011110111010111" => color_data <= "000000000000";
      when "011110111011000" => color_data <= "000000000000";
      when "011110111011001" => color_data <= "000000000000";
      when "011110111011010" => color_data <= "000000000000";
      when "011110111011011" => color_data <= "000000000000";
      when "011110111011100" => color_data <= "000000000000";
      when "011110111011101" => color_data <= "000000000000";
      when "011110111011110" => color_data <= "000000000000";
      when "011110111011111" => color_data <= "000000000000";
      when "011110111100000" => color_data <= "000000000000";
      when "011110111100001" => color_data <= "000000000000";
      when "011110111100010" => color_data <= "000000000000";
      when "011110111100011" => color_data <= "000000000000";
      when "011111000000000" => color_data <= "000000000000";
      when "011111000000001" => color_data <= "000000000000";
      when "011111000000010" => color_data <= "000000000000";
      when "011111000000011" => color_data <= "000000000000";
      when "011111000000100" => color_data <= "000000000000";
      when "011111000000101" => color_data <= "000000000000";
      when "011111000000110" => color_data <= "000000000000";
      when "011111000000111" => color_data <= "000000000000";
      when "011111000001000" => color_data <= "000000000000";
      when "011111000001001" => color_data <= "000000000000";
      when "011111000001010" => color_data <= "000000000000";
      when "011111000001011" => color_data <= "000000000000";
      when "011111000001100" => color_data <= "000000000000";
      when "011111000001101" => color_data <= "000000000000";
      when "011111000001110" => color_data <= "000000000000";
      when "011111000001111" => color_data <= "000000000000";
      when "011111000010000" => color_data <= "000000000000";
      when "011111000010001" => color_data <= "000000000000";
      when "011111000010010" => color_data <= "000000000000";
      when "011111000010011" => color_data <= "000000000000";
      when "011111000010100" => color_data <= "000000000000";
      when "011111000010101" => color_data <= "000000000000";
      when "011111000010110" => color_data <= "000000000000";
      when "011111000010111" => color_data <= "000000000000";
      when "011111000011000" => color_data <= "000000000000";
      when "011111000011001" => color_data <= "000000000000";
      when "011111000011010" => color_data <= "000000000000";
      when "011111000011011" => color_data <= "000000000000";
      when "011111000011100" => color_data <= "000000000000";
      when "011111000011101" => color_data <= "000000000000";
      when "011111000011110" => color_data <= "000000000000";
      when "011111000011111" => color_data <= "000000000000";
      when "011111000100000" => color_data <= "000000000000";
      when "011111000100001" => color_data <= "010101010011";
      when "011111000100010" => color_data <= "111110110000";
      when "011111000100011" => color_data <= "111111000000";
      when "011111000100100" => color_data <= "111111000000";
      when "011111000100101" => color_data <= "111111000001";
      when "011111000100110" => color_data <= "111111000001";
      when "011111000100111" => color_data <= "111111000001";
      when "011111000101000" => color_data <= "111111000001";
      when "011111000101001" => color_data <= "111111000001";
      when "011111000101010" => color_data <= "111111000001";
      when "011111000101011" => color_data <= "111111000001";
      when "011111000101100" => color_data <= "111111000001";
      when "011111000101101" => color_data <= "111111000001";
      when "011111000101110" => color_data <= "111111000001";
      when "011111000101111" => color_data <= "111111000001";
      when "011111000110000" => color_data <= "111111000001";
      when "011111000110001" => color_data <= "111111000001";
      when "011111000110010" => color_data <= "111111000001";
      when "011111000110011" => color_data <= "111111000001";
      when "011111000110100" => color_data <= "111111000001";
      when "011111000110101" => color_data <= "111111000001";
      when "011111000110110" => color_data <= "111111000001";
      when "011111000110111" => color_data <= "111111000001";
      when "011111000111000" => color_data <= "111111000001";
      when "011111000111001" => color_data <= "111111000001";
      when "011111000111010" => color_data <= "111111000001";
      when "011111000111011" => color_data <= "111111000001";
      when "011111000111100" => color_data <= "111111000001";
      when "011111000111101" => color_data <= "111111000001";
      when "011111000111110" => color_data <= "111111000001";
      when "011111000111111" => color_data <= "111111000001";
      when "011111001000000" => color_data <= "111111000001";
      when "011111001000001" => color_data <= "111111000000";
      when "011111001000010" => color_data <= "111110110000";
      when "011111001000011" => color_data <= "100001110010";
      when "011111001000100" => color_data <= "000000000000";
      when "011111001000101" => color_data <= "000000000000";
      when "011111001000110" => color_data <= "000000000000";
      when "011111001000111" => color_data <= "000000000000";
      when "011111001001000" => color_data <= "000000000000";
      when "011111001001001" => color_data <= "000000000000";
      when "011111001001010" => color_data <= "000000000000";
      when "011111001001011" => color_data <= "000000000000";
      when "011111001001100" => color_data <= "000000000000";
      when "011111001001101" => color_data <= "000000000000";
      when "011111001001110" => color_data <= "000000000000";
      when "011111001001111" => color_data <= "000000000000";
      when "011111001010000" => color_data <= "000000000000";
      when "011111001010001" => color_data <= "000000000000";
      when "011111001010010" => color_data <= "000000000000";
      when "011111001010011" => color_data <= "000000000000";
      when "011111001010100" => color_data <= "000000000000";
      when "011111001010101" => color_data <= "000000000000";
      when "011111001010110" => color_data <= "000000000000";
      when "011111001010111" => color_data <= "000000000000";
      when "011111001011000" => color_data <= "000000000000";
      when "011111001011001" => color_data <= "000000000000";
      when "011111001011010" => color_data <= "000000000000";
      when "011111001011011" => color_data <= "000000000000";
      when "011111001011100" => color_data <= "000000000000";
      when "011111001011101" => color_data <= "000000000000";
      when "011111001011110" => color_data <= "000000000000";
      when "011111001011111" => color_data <= "000000000000";
      when "011111001100000" => color_data <= "000000000000";
      when "011111001100001" => color_data <= "000000000000";
      when "011111001100010" => color_data <= "000000000000";
      when "011111001100011" => color_data <= "000000000000";
      when "011111010000000" => color_data <= "000000000000";
      when "011111010000001" => color_data <= "000000000000";
      when "011111010000010" => color_data <= "000000000000";
      when "011111010000011" => color_data <= "000000000000";
      when "011111010000100" => color_data <= "000000000000";
      when "011111010000101" => color_data <= "000000000000";
      when "011111010000110" => color_data <= "000000000000";
      when "011111010000111" => color_data <= "000000000000";
      when "011111010001000" => color_data <= "000000000000";
      when "011111010001001" => color_data <= "000000000000";
      when "011111010001010" => color_data <= "000000000000";
      when "011111010001011" => color_data <= "000000000000";
      when "011111010001100" => color_data <= "000000000000";
      when "011111010001101" => color_data <= "000000000000";
      when "011111010001110" => color_data <= "000000000000";
      when "011111010001111" => color_data <= "000000000000";
      when "011111010010000" => color_data <= "000000000000";
      when "011111010010001" => color_data <= "000000000000";
      when "011111010010010" => color_data <= "000000000000";
      when "011111010010011" => color_data <= "000000000000";
      when "011111010010100" => color_data <= "000000000000";
      when "011111010010101" => color_data <= "000000000000";
      when "011111010010110" => color_data <= "000000000000";
      when "011111010010111" => color_data <= "000000000000";
      when "011111010011000" => color_data <= "000000000000";
      when "011111010011001" => color_data <= "000000000000";
      when "011111010011010" => color_data <= "000000000000";
      when "011111010011011" => color_data <= "000000000000";
      when "011111010011100" => color_data <= "000000000000";
      when "011111010011101" => color_data <= "000000000000";
      when "011111010011110" => color_data <= "000000000000";
      when "011111010011111" => color_data <= "000000000000";
      when "011111010100000" => color_data <= "000000000000";
      when "011111010100001" => color_data <= "010101000010";
      when "011111010100010" => color_data <= "111111000000";
      when "011111010100011" => color_data <= "111111010001";
      when "011111010100100" => color_data <= "111111010001";
      when "011111010100101" => color_data <= "111111010001";
      when "011111010100110" => color_data <= "111111010001";
      when "011111010100111" => color_data <= "111111010001";
      when "011111010101000" => color_data <= "111111010001";
      when "011111010101001" => color_data <= "111111010001";
      when "011111010101010" => color_data <= "111111010001";
      when "011111010101011" => color_data <= "111111010001";
      when "011111010101100" => color_data <= "111111010001";
      when "011111010101101" => color_data <= "111111010001";
      when "011111010101110" => color_data <= "111111010001";
      when "011111010101111" => color_data <= "111111010001";
      when "011111010110000" => color_data <= "111111010001";
      when "011111010110001" => color_data <= "111111010001";
      when "011111010110010" => color_data <= "111111010001";
      when "011111010110011" => color_data <= "111111010001";
      when "011111010110100" => color_data <= "111111010001";
      when "011111010110101" => color_data <= "111111010001";
      when "011111010110110" => color_data <= "111111010001";
      when "011111010110111" => color_data <= "111111010001";
      when "011111010111000" => color_data <= "111111010001";
      when "011111010111001" => color_data <= "111111010001";
      when "011111010111010" => color_data <= "111111010001";
      when "011111010111011" => color_data <= "111111010001";
      when "011111010111100" => color_data <= "111111010001";
      when "011111010111101" => color_data <= "111111010001";
      when "011111010111110" => color_data <= "111111010001";
      when "011111010111111" => color_data <= "111111010001";
      when "011111011000000" => color_data <= "111111010001";
      when "011111011000001" => color_data <= "111111010001";
      when "011111011000010" => color_data <= "111111000000";
      when "011111011000011" => color_data <= "100001110011";
      when "011111011000100" => color_data <= "000000000000";
      when "011111011000101" => color_data <= "000000000000";
      when "011111011000110" => color_data <= "000000000000";
      when "011111011000111" => color_data <= "000000000000";
      when "011111011001000" => color_data <= "000000000000";
      when "011111011001001" => color_data <= "000000000000";
      when "011111011001010" => color_data <= "000000000000";
      when "011111011001011" => color_data <= "000000000000";
      when "011111011001100" => color_data <= "000000000000";
      when "011111011001101" => color_data <= "000000000000";
      when "011111011001110" => color_data <= "000000000000";
      when "011111011001111" => color_data <= "000000000000";
      when "011111011010000" => color_data <= "000000000000";
      when "011111011010001" => color_data <= "000000000000";
      when "011111011010010" => color_data <= "000000000000";
      when "011111011010011" => color_data <= "000000000000";
      when "011111011010100" => color_data <= "000000000000";
      when "011111011010101" => color_data <= "000000000000";
      when "011111011010110" => color_data <= "000000000000";
      when "011111011010111" => color_data <= "000000000000";
      when "011111011011000" => color_data <= "000000000000";
      when "011111011011001" => color_data <= "000000000000";
      when "011111011011010" => color_data <= "000000000000";
      when "011111011011011" => color_data <= "000000000000";
      when "011111011011100" => color_data <= "000000000000";
      when "011111011011101" => color_data <= "000000000000";
      when "011111011011110" => color_data <= "000000000000";
      when "011111011011111" => color_data <= "000000000000";
      when "011111011100000" => color_data <= "000000000000";
      when "011111011100001" => color_data <= "000000000000";
      when "011111011100010" => color_data <= "000000000000";
      when "011111011100011" => color_data <= "000000000000";
      when "011111100000000" => color_data <= "000000000000";
      when "011111100000001" => color_data <= "000000000000";
      when "011111100000010" => color_data <= "000000000000";
      when "011111100000011" => color_data <= "000000000000";
      when "011111100000100" => color_data <= "000000000000";
      when "011111100000101" => color_data <= "000000000000";
      when "011111100000110" => color_data <= "000000000000";
      when "011111100000111" => color_data <= "000000000000";
      when "011111100001000" => color_data <= "000000000000";
      when "011111100001001" => color_data <= "000000000000";
      when "011111100001010" => color_data <= "000000000000";
      when "011111100001011" => color_data <= "000000000000";
      when "011111100001100" => color_data <= "000000000000";
      when "011111100001101" => color_data <= "000000000000";
      when "011111100001110" => color_data <= "000000000000";
      when "011111100001111" => color_data <= "000000000000";
      when "011111100010000" => color_data <= "000000000000";
      when "011111100010001" => color_data <= "000000000000";
      when "011111100010010" => color_data <= "000000000000";
      when "011111100010011" => color_data <= "000000000000";
      when "011111100010100" => color_data <= "000000000000";
      when "011111100010101" => color_data <= "000000000000";
      when "011111100010110" => color_data <= "000000000000";
      when "011111100010111" => color_data <= "000000000000";
      when "011111100011000" => color_data <= "000000000000";
      when "011111100011001" => color_data <= "000000000000";
      when "011111100011010" => color_data <= "000000000000";
      when "011111100011011" => color_data <= "000000000000";
      when "011111100011100" => color_data <= "000000000000";
      when "011111100011101" => color_data <= "000000000000";
      when "011111100011110" => color_data <= "000000000000";
      when "011111100011111" => color_data <= "000000000000";
      when "011111100100000" => color_data <= "000000000000";
      when "011111100100001" => color_data <= "010101000011";
      when "011111100100010" => color_data <= "110110010000";
      when "011111100100011" => color_data <= "111010100001";
      when "011111100100100" => color_data <= "111010100001";
      when "011111100100101" => color_data <= "111010100001";
      when "011111100100110" => color_data <= "111010100001";
      when "011111100100111" => color_data <= "111010100001";
      when "011111100101000" => color_data <= "111010100001";
      when "011111100101001" => color_data <= "111010100001";
      when "011111100101010" => color_data <= "111010100001";
      when "011111100101011" => color_data <= "111010100001";
      when "011111100101100" => color_data <= "111010100001";
      when "011111100101101" => color_data <= "111010100001";
      when "011111100101110" => color_data <= "111010100001";
      when "011111100101111" => color_data <= "111010100001";
      when "011111100110000" => color_data <= "111010100001";
      when "011111100110001" => color_data <= "111010100001";
      when "011111100110010" => color_data <= "111010100001";
      when "011111100110011" => color_data <= "111010100001";
      when "011111100110100" => color_data <= "111010100001";
      when "011111100110101" => color_data <= "111010100001";
      when "011111100110110" => color_data <= "111010100001";
      when "011111100110111" => color_data <= "111010100001";
      when "011111100111000" => color_data <= "111010100001";
      when "011111100111001" => color_data <= "111010100001";
      when "011111100111010" => color_data <= "111010100001";
      when "011111100111011" => color_data <= "111010100001";
      when "011111100111100" => color_data <= "111010100001";
      when "011111100111101" => color_data <= "111010100001";
      when "011111100111110" => color_data <= "111010100001";
      when "011111100111111" => color_data <= "111010100001";
      when "011111101000000" => color_data <= "111010100001";
      when "011111101000001" => color_data <= "111010100001";
      when "011111101000010" => color_data <= "111010100000";
      when "011111101000011" => color_data <= "011101100010";
      when "011111101000100" => color_data <= "000100010001";
      when "011111101000101" => color_data <= "000000000000";
      when "011111101000110" => color_data <= "000000000000";
      when "011111101000111" => color_data <= "000000000000";
      when "011111101001000" => color_data <= "000000000000";
      when "011111101001001" => color_data <= "000000000000";
      when "011111101001010" => color_data <= "000000000000";
      when "011111101001011" => color_data <= "000000000000";
      when "011111101001100" => color_data <= "000000000000";
      when "011111101001101" => color_data <= "000000000000";
      when "011111101001110" => color_data <= "000000000000";
      when "011111101001111" => color_data <= "000000000000";
      when "011111101010000" => color_data <= "000000000000";
      when "011111101010001" => color_data <= "000000000000";
      when "011111101010010" => color_data <= "000000000000";
      when "011111101010011" => color_data <= "000000000000";
      when "011111101010100" => color_data <= "000000000000";
      when "011111101010101" => color_data <= "000000000000";
      when "011111101010110" => color_data <= "000000000000";
      when "011111101010111" => color_data <= "000000000000";
      when "011111101011000" => color_data <= "000000000000";
      when "011111101011001" => color_data <= "000000000000";
      when "011111101011010" => color_data <= "000000000000";
      when "011111101011011" => color_data <= "000000000000";
      when "011111101011100" => color_data <= "000000000000";
      when "011111101011101" => color_data <= "000000000000";
      when "011111101011110" => color_data <= "000000000000";
      when "011111101011111" => color_data <= "000000000000";
      when "011111101100000" => color_data <= "000000000000";
      when "011111101100001" => color_data <= "000000000000";
      when "011111101100010" => color_data <= "000000000000";
      when "011111101100011" => color_data <= "000000000000";
      when "011111110000000" => color_data <= "000000000000";
      when "011111110000001" => color_data <= "000000000000";
      when "011111110000010" => color_data <= "000000000000";
      when "011111110000011" => color_data <= "000000000000";
      when "011111110000100" => color_data <= "000000000000";
      when "011111110000101" => color_data <= "000000000000";
      when "011111110000110" => color_data <= "000000000000";
      when "011111110000111" => color_data <= "000000000000";
      when "011111110001000" => color_data <= "000000000000";
      when "011111110001001" => color_data <= "000000000000";
      when "011111110001010" => color_data <= "000000000000";
      when "011111110001011" => color_data <= "000000000000";
      when "011111110001100" => color_data <= "000000000000";
      when "011111110001101" => color_data <= "000000000000";
      when "011111110001110" => color_data <= "000000000000";
      when "011111110001111" => color_data <= "000000000000";
      when "011111110010000" => color_data <= "000000000000";
      when "011111110010001" => color_data <= "000000000000";
      when "011111110010010" => color_data <= "000000000000";
      when "011111110010011" => color_data <= "000000000000";
      when "011111110010100" => color_data <= "000000000000";
      when "011111110010101" => color_data <= "000000000000";
      when "011111110010110" => color_data <= "000000000000";
      when "011111110010111" => color_data <= "000000000000";
      when "011111110011000" => color_data <= "000000000000";
      when "011111110011001" => color_data <= "000000000000";
      when "011111110011010" => color_data <= "000000000000";
      when "011111110011011" => color_data <= "000000000000";
      when "011111110011100" => color_data <= "000000000000";
      when "011111110011101" => color_data <= "000000000000";
      when "011111110011110" => color_data <= "000000000000";
      when "011111110011111" => color_data <= "000100010001";
      when "011111110100000" => color_data <= "010000110010";
      when "011111110100001" => color_data <= "010100110010";
      when "011111110100010" => color_data <= "011000110001";
      when "011111110100011" => color_data <= "011000110010";
      when "011111110100100" => color_data <= "011000110010";
      when "011111110100101" => color_data <= "011000110010";
      when "011111110100110" => color_data <= "011000110010";
      when "011111110100111" => color_data <= "011000110010";
      when "011111110101000" => color_data <= "011000110010";
      when "011111110101001" => color_data <= "011000110010";
      when "011111110101010" => color_data <= "011000110010";
      when "011111110101011" => color_data <= "011000110010";
      when "011111110101100" => color_data <= "011000110010";
      when "011111110101101" => color_data <= "011000110010";
      when "011111110101110" => color_data <= "011000110010";
      when "011111110101111" => color_data <= "011000110010";
      when "011111110110000" => color_data <= "011000110010";
      when "011111110110001" => color_data <= "011000110010";
      when "011111110110010" => color_data <= "011000110010";
      when "011111110110011" => color_data <= "011000110010";
      when "011111110110100" => color_data <= "011000110010";
      when "011111110110101" => color_data <= "011000110010";
      when "011111110110110" => color_data <= "011000110010";
      when "011111110110111" => color_data <= "011000110010";
      when "011111110111000" => color_data <= "011000110010";
      when "011111110111001" => color_data <= "011000110010";
      when "011111110111010" => color_data <= "011000110010";
      when "011111110111011" => color_data <= "011000110010";
      when "011111110111100" => color_data <= "011000110010";
      when "011111110111101" => color_data <= "011000110010";
      when "011111110111110" => color_data <= "011000110010";
      when "011111110111111" => color_data <= "011000110010";
      when "011111111000000" => color_data <= "011000110010";
      when "011111111000001" => color_data <= "011000110010";
      when "011111111000010" => color_data <= "011100110010";
      when "011111111000011" => color_data <= "011000110010";
      when "011111111000100" => color_data <= "010000010000";
      when "011111111000101" => color_data <= "010000110011";
      when "011111111000110" => color_data <= "000000000000";
      when "011111111000111" => color_data <= "000000000000";
      when "011111111001000" => color_data <= "000000000000";
      when "011111111001001" => color_data <= "000000000000";
      when "011111111001010" => color_data <= "000000000000";
      when "011111111001011" => color_data <= "000000000000";
      when "011111111001100" => color_data <= "000000000000";
      when "011111111001101" => color_data <= "000000000000";
      when "011111111001110" => color_data <= "000000000000";
      when "011111111001111" => color_data <= "000000000000";
      when "011111111010000" => color_data <= "000000000000";
      when "011111111010001" => color_data <= "000000000000";
      when "011111111010010" => color_data <= "000000000000";
      when "011111111010011" => color_data <= "000000000000";
      when "011111111010100" => color_data <= "000000000000";
      when "011111111010101" => color_data <= "000000000000";
      when "011111111010110" => color_data <= "000000000000";
      when "011111111010111" => color_data <= "000000000000";
      when "011111111011000" => color_data <= "000000000000";
      when "011111111011001" => color_data <= "000000000000";
      when "011111111011010" => color_data <= "000000000000";
      when "011111111011011" => color_data <= "000000000000";
      when "011111111011100" => color_data <= "000000000000";
      when "011111111011101" => color_data <= "000000000000";
      when "011111111011110" => color_data <= "000000000000";
      when "011111111011111" => color_data <= "000000000000";
      when "011111111100000" => color_data <= "000000000000";
      when "011111111100001" => color_data <= "000000000000";
      when "011111111100010" => color_data <= "000000000000";
      when "011111111100011" => color_data <= "000000000000";
      when "100000000000000" => color_data <= "000000000000";
      when "100000000000001" => color_data <= "000000000000";
      when "100000000000010" => color_data <= "000000000000";
      when "100000000000011" => color_data <= "000000000000";
      when "100000000000100" => color_data <= "000000000000";
      when "100000000000101" => color_data <= "000000000000";
      when "100000000000110" => color_data <= "000000000000";
      when "100000000000111" => color_data <= "000000000000";
      when "100000000001000" => color_data <= "000000000000";
      when "100000000001001" => color_data <= "000000000000";
      when "100000000001010" => color_data <= "000000000000";
      when "100000000001011" => color_data <= "000000000000";
      when "100000000001100" => color_data <= "000000000000";
      when "100000000001101" => color_data <= "000000000000";
      when "100000000001110" => color_data <= "000000000000";
      when "100000000001111" => color_data <= "000000000000";
      when "100000000010000" => color_data <= "000000000000";
      when "100000000010001" => color_data <= "000000000000";
      when "100000000010010" => color_data <= "000000000000";
      when "100000000010011" => color_data <= "000000000000";
      when "100000000010100" => color_data <= "000000000000";
      when "100000000010101" => color_data <= "000000000000";
      when "100000000010110" => color_data <= "000000000000";
      when "100000000010111" => color_data <= "000000000000";
      when "100000000011000" => color_data <= "000000000000";
      when "100000000011001" => color_data <= "000000000000";
      when "100000000011010" => color_data <= "000000000000";
      when "100000000011011" => color_data <= "000000000000";
      when "100000000011100" => color_data <= "000000000000";
      when "100000000011101" => color_data <= "000000000000";
      when "100000000011110" => color_data <= "000000000000";
      when "100000000011111" => color_data <= "001000100010";
      when "100000000100000" => color_data <= "010100010000";
      when "100000000100001" => color_data <= "011100110001";
      when "100000000100010" => color_data <= "011101000010";
      when "100000000100011" => color_data <= "011101000001";
      when "100000000100100" => color_data <= "011101000001";
      when "100000000100101" => color_data <= "011101000001";
      when "100000000100110" => color_data <= "011101000010";
      when "100000000100111" => color_data <= "011101000010";
      when "100000000101000" => color_data <= "011101000010";
      when "100000000101001" => color_data <= "011101000010";
      when "100000000101010" => color_data <= "011101000010";
      when "100000000101011" => color_data <= "011101000010";
      when "100000000101100" => color_data <= "011101000010";
      when "100000000101101" => color_data <= "011101000010";
      when "100000000101110" => color_data <= "011101000010";
      when "100000000101111" => color_data <= "011101000010";
      when "100000000110000" => color_data <= "011101000010";
      when "100000000110001" => color_data <= "011101000010";
      when "100000000110010" => color_data <= "011101000010";
      when "100000000110011" => color_data <= "011101000010";
      when "100000000110100" => color_data <= "011101000010";
      when "100000000110101" => color_data <= "011101000010";
      when "100000000110110" => color_data <= "011101000010";
      when "100000000110111" => color_data <= "011101000010";
      when "100000000111000" => color_data <= "011101000010";
      when "100000000111001" => color_data <= "011101000010";
      when "100000000111010" => color_data <= "011101000010";
      when "100000000111011" => color_data <= "011101000010";
      when "100000000111100" => color_data <= "011101000010";
      when "100000000111101" => color_data <= "011101000010";
      when "100000000111110" => color_data <= "011101000010";
      when "100000000111111" => color_data <= "011101000010";
      when "100000001000000" => color_data <= "011101000010";
      when "100000001000001" => color_data <= "011101000001";
      when "100000001000010" => color_data <= "011101000010";
      when "100000001000011" => color_data <= "011101000001";
      when "100000001000100" => color_data <= "010100010000";
      when "100000001000101" => color_data <= "010000110011";
      when "100000001000110" => color_data <= "000000000000";
      when "100000001000111" => color_data <= "000000000000";
      when "100000001001000" => color_data <= "000000000000";
      when "100000001001001" => color_data <= "000000000000";
      when "100000001001010" => color_data <= "000000000000";
      when "100000001001011" => color_data <= "000000000000";
      when "100000001001100" => color_data <= "000000000000";
      when "100000001001101" => color_data <= "000000000000";
      when "100000001001110" => color_data <= "000000000000";
      when "100000001001111" => color_data <= "000000000000";
      when "100000001010000" => color_data <= "000000000000";
      when "100000001010001" => color_data <= "000000000000";
      when "100000001010010" => color_data <= "000000000000";
      when "100000001010011" => color_data <= "000000000000";
      when "100000001010100" => color_data <= "000000000000";
      when "100000001010101" => color_data <= "000000000000";
      when "100000001010110" => color_data <= "000000000000";
      when "100000001010111" => color_data <= "000000000000";
      when "100000001011000" => color_data <= "000000000000";
      when "100000001011001" => color_data <= "000000000000";
      when "100000001011010" => color_data <= "000000000000";
      when "100000001011011" => color_data <= "000000000000";
      when "100000001011100" => color_data <= "000000000000";
      when "100000001011101" => color_data <= "000000000000";
      when "100000001011110" => color_data <= "000000000000";
      when "100000001011111" => color_data <= "000000000000";
      when "100000001100000" => color_data <= "000000000000";
      when "100000001100001" => color_data <= "000000000000";
      when "100000001100010" => color_data <= "000000000000";
      when "100000001100011" => color_data <= "000000000000";
      when "100000010000000" => color_data <= "000000000000";
      when "100000010000001" => color_data <= "000000000000";
      when "100000010000010" => color_data <= "000000000000";
      when "100000010000011" => color_data <= "000000000000";
      when "100000010000100" => color_data <= "000000000000";
      when "100000010000101" => color_data <= "000000000000";
      when "100000010000110" => color_data <= "000000000000";
      when "100000010000111" => color_data <= "000000000000";
      when "100000010001000" => color_data <= "000000000000";
      when "100000010001001" => color_data <= "000000000000";
      when "100000010001010" => color_data <= "000000000000";
      when "100000010001011" => color_data <= "000000000000";
      when "100000010001100" => color_data <= "000000000000";
      when "100000010001101" => color_data <= "000000000000";
      when "100000010001110" => color_data <= "000000000000";
      when "100000010001111" => color_data <= "000000000000";
      when "100000010010000" => color_data <= "000000000000";
      when "100000010010001" => color_data <= "000000000000";
      when "100000010010010" => color_data <= "000000000000";
      when "100000010010011" => color_data <= "000000000000";
      when "100000010010100" => color_data <= "000000000000";
      when "100000010010101" => color_data <= "000000000000";
      when "100000010010110" => color_data <= "000000000000";
      when "100000010010111" => color_data <= "000000000000";
      when "100000010011000" => color_data <= "000000000000";
      when "100000010011001" => color_data <= "000000000000";
      when "100000010011010" => color_data <= "000000000000";
      when "100000010011011" => color_data <= "000000000000";
      when "100000010011100" => color_data <= "000000000000";
      when "100000010011101" => color_data <= "000000000000";
      when "100000010011110" => color_data <= "000000000000";
      when "100000010011111" => color_data <= "001000100010";
      when "100000010100000" => color_data <= "011000100000";
      when "100000010100001" => color_data <= "011101000010";
      when "100000010100010" => color_data <= "011101000010";
      when "100000010100011" => color_data <= "011101000010";
      when "100000010100100" => color_data <= "011101000010";
      when "100000010100101" => color_data <= "011101000010";
      when "100000010100110" => color_data <= "011101000010";
      when "100000010100111" => color_data <= "011101000010";
      when "100000010101000" => color_data <= "011101000010";
      when "100000010101001" => color_data <= "011101000010";
      when "100000010101010" => color_data <= "011101000010";
      when "100000010101011" => color_data <= "011101000010";
      when "100000010101100" => color_data <= "011101000010";
      when "100000010101101" => color_data <= "011101000010";
      when "100000010101110" => color_data <= "011101000010";
      when "100000010101111" => color_data <= "011101000010";
      when "100000010110000" => color_data <= "011101000010";
      when "100000010110001" => color_data <= "011101000010";
      when "100000010110010" => color_data <= "011101000010";
      when "100000010110011" => color_data <= "011101000010";
      when "100000010110100" => color_data <= "011101000010";
      when "100000010110101" => color_data <= "011101000010";
      when "100000010110110" => color_data <= "011101000010";
      when "100000010110111" => color_data <= "011101000010";
      when "100000010111000" => color_data <= "011101000010";
      when "100000010111001" => color_data <= "011101000010";
      when "100000010111010" => color_data <= "011101000010";
      when "100000010111011" => color_data <= "011101000010";
      when "100000010111100" => color_data <= "011101000010";
      when "100000010111101" => color_data <= "011101000010";
      when "100000010111110" => color_data <= "011101000010";
      when "100000010111111" => color_data <= "011101000010";
      when "100000011000000" => color_data <= "011101000010";
      when "100000011000001" => color_data <= "011101000010";
      when "100000011000010" => color_data <= "011101000010";
      when "100000011000011" => color_data <= "011101000010";
      when "100000011000100" => color_data <= "010100100000";
      when "100000011000101" => color_data <= "010000110011";
      when "100000011000110" => color_data <= "000000000000";
      when "100000011000111" => color_data <= "000000000000";
      when "100000011001000" => color_data <= "000000000000";
      when "100000011001001" => color_data <= "000000000000";
      when "100000011001010" => color_data <= "000000000000";
      when "100000011001011" => color_data <= "000000000000";
      when "100000011001100" => color_data <= "000000000000";
      when "100000011001101" => color_data <= "000000000000";
      when "100000011001110" => color_data <= "000000000000";
      when "100000011001111" => color_data <= "000000000000";
      when "100000011010000" => color_data <= "000000000000";
      when "100000011010001" => color_data <= "000000000000";
      when "100000011010010" => color_data <= "000000000000";
      when "100000011010011" => color_data <= "000000000000";
      when "100000011010100" => color_data <= "000000000000";
      when "100000011010101" => color_data <= "000000000000";
      when "100000011010110" => color_data <= "000000000000";
      when "100000011010111" => color_data <= "000000000000";
      when "100000011011000" => color_data <= "000000000000";
      when "100000011011001" => color_data <= "000000000000";
      when "100000011011010" => color_data <= "000000000000";
      when "100000011011011" => color_data <= "000000000000";
      when "100000011011100" => color_data <= "000000000000";
      when "100000011011101" => color_data <= "000000000000";
      when "100000011011110" => color_data <= "000000000000";
      when "100000011011111" => color_data <= "000000000000";
      when "100000011100000" => color_data <= "000000000000";
      when "100000011100001" => color_data <= "000000000000";
      when "100000011100010" => color_data <= "000000000000";
      when "100000011100011" => color_data <= "000000000000";
      when "100000100000000" => color_data <= "000000000000";
      when "100000100000001" => color_data <= "000000000000";
      when "100000100000010" => color_data <= "000000000000";
      when "100000100000011" => color_data <= "000000000000";
      when "100000100000100" => color_data <= "000000000000";
      when "100000100000101" => color_data <= "000000000000";
      when "100000100000110" => color_data <= "000000000000";
      when "100000100000111" => color_data <= "000000000000";
      when "100000100001000" => color_data <= "000000000000";
      when "100000100001001" => color_data <= "000000000000";
      when "100000100001010" => color_data <= "000000000000";
      when "100000100001011" => color_data <= "000000000000";
      when "100000100001100" => color_data <= "000000000000";
      when "100000100001101" => color_data <= "000000000000";
      when "100000100001110" => color_data <= "000000000000";
      when "100000100001111" => color_data <= "000000000000";
      when "100000100010000" => color_data <= "000000000000";
      when "100000100010001" => color_data <= "000000000000";
      when "100000100010010" => color_data <= "000000000000";
      when "100000100010011" => color_data <= "000000000000";
      when "100000100010100" => color_data <= "000000000000";
      when "100000100010101" => color_data <= "000000000000";
      when "100000100010110" => color_data <= "000000000000";
      when "100000100010111" => color_data <= "000000000000";
      when "100000100011000" => color_data <= "000000000000";
      when "100000100011001" => color_data <= "000000000000";
      when "100000100011010" => color_data <= "000000000000";
      when "100000100011011" => color_data <= "000000000000";
      when "100000100011100" => color_data <= "000000000000";
      when "100000100011101" => color_data <= "000000000000";
      when "100000100011110" => color_data <= "000000000000";
      when "100000100011111" => color_data <= "000100010001";
      when "100000100100000" => color_data <= "010100100000";
      when "100000100100001" => color_data <= "011101000010";
      when "100000100100010" => color_data <= "011101000010";
      when "100000100100011" => color_data <= "011101000010";
      when "100000100100100" => color_data <= "011101000010";
      when "100000100100101" => color_data <= "011101000010";
      when "100000100100110" => color_data <= "011101000010";
      when "100000100100111" => color_data <= "011101000010";
      when "100000100101000" => color_data <= "011101000010";
      when "100000100101001" => color_data <= "011101000010";
      when "100000100101010" => color_data <= "011101000010";
      when "100000100101011" => color_data <= "011101000010";
      when "100000100101100" => color_data <= "011101000010";
      when "100000100101101" => color_data <= "011101000010";
      when "100000100101110" => color_data <= "011101000010";
      when "100000100101111" => color_data <= "011101000010";
      when "100000100110000" => color_data <= "011101000010";
      when "100000100110001" => color_data <= "011101000010";
      when "100000100110010" => color_data <= "011101000010";
      when "100000100110011" => color_data <= "011101000010";
      when "100000100110100" => color_data <= "011101000010";
      when "100000100110101" => color_data <= "011101000010";
      when "100000100110110" => color_data <= "011101000010";
      when "100000100110111" => color_data <= "011101000010";
      when "100000100111000" => color_data <= "011101000010";
      when "100000100111001" => color_data <= "011101000010";
      when "100000100111010" => color_data <= "011101000010";
      when "100000100111011" => color_data <= "011101000010";
      when "100000100111100" => color_data <= "011101000010";
      when "100000100111101" => color_data <= "011101000010";
      when "100000100111110" => color_data <= "011101000010";
      when "100000100111111" => color_data <= "011101000010";
      when "100000101000000" => color_data <= "011101000010";
      when "100000101000001" => color_data <= "011101000010";
      when "100000101000010" => color_data <= "011101000010";
      when "100000101000011" => color_data <= "011101000010";
      when "100000101000100" => color_data <= "010100010000";
      when "100000101000101" => color_data <= "010000110010";
      when "100000101000110" => color_data <= "000000000000";
      when "100000101000111" => color_data <= "000000000000";
      when "100000101001000" => color_data <= "000000000000";
      when "100000101001001" => color_data <= "000000000000";
      when "100000101001010" => color_data <= "000000000000";
      when "100000101001011" => color_data <= "000000000000";
      when "100000101001100" => color_data <= "000000000000";
      when "100000101001101" => color_data <= "000000000000";
      when "100000101001110" => color_data <= "000000000000";
      when "100000101001111" => color_data <= "000000000000";
      when "100000101010000" => color_data <= "000000000000";
      when "100000101010001" => color_data <= "000000000000";
      when "100000101010010" => color_data <= "000000000000";
      when "100000101010011" => color_data <= "000000000000";
      when "100000101010100" => color_data <= "000000000000";
      when "100000101010101" => color_data <= "000000000000";
      when "100000101010110" => color_data <= "000000000000";
      when "100000101010111" => color_data <= "000000000000";
      when "100000101011000" => color_data <= "000000000000";
      when "100000101011001" => color_data <= "000000000000";
      when "100000101011010" => color_data <= "000000000000";
      when "100000101011011" => color_data <= "000000000000";
      when "100000101011100" => color_data <= "000000000000";
      when "100000101011101" => color_data <= "000000000000";
      when "100000101011110" => color_data <= "000000000000";
      when "100000101011111" => color_data <= "000000000000";
      when "100000101100000" => color_data <= "000000000000";
      when "100000101100001" => color_data <= "000000000000";
      when "100000101100010" => color_data <= "000000000000";
      when "100000101100011" => color_data <= "000000000000";
      when "100000110000000" => color_data <= "000000000000";
      when "100000110000001" => color_data <= "000000000000";
      when "100000110000010" => color_data <= "000000000000";
      when "100000110000011" => color_data <= "000000000000";
      when "100000110000100" => color_data <= "000000000000";
      when "100000110000101" => color_data <= "000000000000";
      when "100000110000110" => color_data <= "000000000000";
      when "100000110000111" => color_data <= "000000000000";
      when "100000110001000" => color_data <= "000000000000";
      when "100000110001001" => color_data <= "000000000000";
      when "100000110001010" => color_data <= "000000000000";
      when "100000110001011" => color_data <= "000000000000";
      when "100000110001100" => color_data <= "000000000000";
      when "100000110001101" => color_data <= "000000000000";
      when "100000110001110" => color_data <= "000000000000";
      when "100000110001111" => color_data <= "000000000000";
      when "100000110010000" => color_data <= "000000000000";
      when "100000110010001" => color_data <= "000000000000";
      when "100000110010010" => color_data <= "000000000000";
      when "100000110010011" => color_data <= "000000000000";
      when "100000110010100" => color_data <= "000000000000";
      when "100000110010101" => color_data <= "000000000000";
      when "100000110010110" => color_data <= "000000000000";
      when "100000110010111" => color_data <= "000000000000";
      when "100000110011000" => color_data <= "000000000000";
      when "100000110011001" => color_data <= "000000000000";
      when "100000110011010" => color_data <= "000000000000";
      when "100000110011011" => color_data <= "000100000000";
      when "100000110011100" => color_data <= "001000100010";
      when "100000110011101" => color_data <= "001000100010";
      when "100000110011110" => color_data <= "001000100001";
      when "100000110011111" => color_data <= "010000110011";
      when "100000110100000" => color_data <= "011000110000";
      when "100000110100001" => color_data <= "011101000010";
      when "100000110100010" => color_data <= "011101000010";
      when "100000110100011" => color_data <= "011101000010";
      when "100000110100100" => color_data <= "011101000010";
      when "100000110100101" => color_data <= "011101000010";
      when "100000110100110" => color_data <= "011101000010";
      when "100000110100111" => color_data <= "011101000010";
      when "100000110101000" => color_data <= "011101000010";
      when "100000110101001" => color_data <= "011101000010";
      when "100000110101010" => color_data <= "011101000010";
      when "100000110101011" => color_data <= "011101000010";
      when "100000110101100" => color_data <= "011101000010";
      when "100000110101101" => color_data <= "011101000010";
      when "100000110101110" => color_data <= "011101000010";
      when "100000110101111" => color_data <= "011101000010";
      when "100000110110000" => color_data <= "011101000010";
      when "100000110110001" => color_data <= "011101000010";
      when "100000110110010" => color_data <= "011101000010";
      when "100000110110011" => color_data <= "011101000010";
      when "100000110110100" => color_data <= "011101000010";
      when "100000110110101" => color_data <= "011101000010";
      when "100000110110110" => color_data <= "011101000010";
      when "100000110110111" => color_data <= "011101000010";
      when "100000110111000" => color_data <= "011101000010";
      when "100000110111001" => color_data <= "011101000010";
      when "100000110111010" => color_data <= "011101000010";
      when "100000110111011" => color_data <= "011101000010";
      when "100000110111100" => color_data <= "011101000010";
      when "100000110111101" => color_data <= "011101000010";
      when "100000110111110" => color_data <= "011101000010";
      when "100000110111111" => color_data <= "011101000010";
      when "100000111000000" => color_data <= "011101000010";
      when "100000111000001" => color_data <= "011101000010";
      when "100000111000010" => color_data <= "011101000010";
      when "100000111000011" => color_data <= "011101000010";
      when "100000111000100" => color_data <= "011000110000";
      when "100000111000101" => color_data <= "010000110010";
      when "100000111000110" => color_data <= "001000100001";
      when "100000111000111" => color_data <= "001000100010";
      when "100000111001000" => color_data <= "001000100010";
      when "100000111001001" => color_data <= "001000100010";
      when "100000111001010" => color_data <= "001000100010";
      when "100000111001011" => color_data <= "000000000000";
      when "100000111001100" => color_data <= "000000000000";
      when "100000111001101" => color_data <= "000000000000";
      when "100000111001110" => color_data <= "000000000000";
      when "100000111001111" => color_data <= "000000000000";
      when "100000111010000" => color_data <= "000000000000";
      when "100000111010001" => color_data <= "000000000000";
      when "100000111010010" => color_data <= "000000000000";
      when "100000111010011" => color_data <= "000000000000";
      when "100000111010100" => color_data <= "000000000000";
      when "100000111010101" => color_data <= "000000000000";
      when "100000111010110" => color_data <= "000000000000";
      when "100000111010111" => color_data <= "000000000000";
      when "100000111011000" => color_data <= "000000000000";
      when "100000111011001" => color_data <= "000000000000";
      when "100000111011010" => color_data <= "000000000000";
      when "100000111011011" => color_data <= "000000000000";
      when "100000111011100" => color_data <= "000000000000";
      when "100000111011101" => color_data <= "000000000000";
      when "100000111011110" => color_data <= "000000000000";
      when "100000111011111" => color_data <= "000000000000";
      when "100000111100000" => color_data <= "000000000000";
      when "100000111100001" => color_data <= "000000000000";
      when "100000111100010" => color_data <= "000000000000";
      when "100000111100011" => color_data <= "000000000000";
      when "100001000000000" => color_data <= "000000000000";
      when "100001000000001" => color_data <= "000000000000";
      when "100001000000010" => color_data <= "000000000000";
      when "100001000000011" => color_data <= "000000000000";
      when "100001000000100" => color_data <= "000000000000";
      when "100001000000101" => color_data <= "000000000000";
      when "100001000000110" => color_data <= "000000000000";
      when "100001000000111" => color_data <= "000000000000";
      when "100001000001000" => color_data <= "000000000000";
      when "100001000001001" => color_data <= "000000000000";
      when "100001000001010" => color_data <= "000000000000";
      when "100001000001011" => color_data <= "000000000000";
      when "100001000001100" => color_data <= "000000000000";
      when "100001000001101" => color_data <= "000000000000";
      when "100001000001110" => color_data <= "000000000000";
      when "100001000001111" => color_data <= "000000000000";
      when "100001000010000" => color_data <= "000000000000";
      when "100001000010001" => color_data <= "000000000000";
      when "100001000010010" => color_data <= "000000000000";
      when "100001000010011" => color_data <= "000000000000";
      when "100001000010100" => color_data <= "000000000000";
      when "100001000010101" => color_data <= "000000000000";
      when "100001000010110" => color_data <= "000000000000";
      when "100001000010111" => color_data <= "000000000000";
      when "100001000011000" => color_data <= "000000000000";
      when "100001000011001" => color_data <= "000000000000";
      when "100001000011010" => color_data <= "000000000000";
      when "100001000011011" => color_data <= "010000110011";
      when "100001000011100" => color_data <= "010000000000";
      when "100001000011101" => color_data <= "011000100000";
      when "100001000011110" => color_data <= "011000100000";
      when "100001000011111" => color_data <= "011000110000";
      when "100001000100000" => color_data <= "011101000010";
      when "100001000100001" => color_data <= "011101000001";
      when "100001000100010" => color_data <= "011100110001";
      when "100001000100011" => color_data <= "011100110001";
      when "100001000100100" => color_data <= "011100110001";
      when "100001000100101" => color_data <= "011100110001";
      when "100001000100110" => color_data <= "011100110001";
      when "100001000100111" => color_data <= "011100110001";
      when "100001000101000" => color_data <= "011100110001";
      when "100001000101001" => color_data <= "011100110001";
      when "100001000101010" => color_data <= "011100110001";
      when "100001000101011" => color_data <= "011100110001";
      when "100001000101100" => color_data <= "011100110001";
      when "100001000101101" => color_data <= "011100110001";
      when "100001000101110" => color_data <= "011100110001";
      when "100001000101111" => color_data <= "011100110001";
      when "100001000110000" => color_data <= "011100110001";
      when "100001000110001" => color_data <= "011100110001";
      when "100001000110010" => color_data <= "011100110001";
      when "100001000110011" => color_data <= "011100110001";
      when "100001000110100" => color_data <= "011100110001";
      when "100001000110101" => color_data <= "011100110001";
      when "100001000110110" => color_data <= "011100110001";
      when "100001000110111" => color_data <= "011100110001";
      when "100001000111000" => color_data <= "011100110001";
      when "100001000111001" => color_data <= "011100110001";
      when "100001000111010" => color_data <= "011100110001";
      when "100001000111011" => color_data <= "011100110001";
      when "100001000111100" => color_data <= "011100110001";
      when "100001000111101" => color_data <= "011100110001";
      when "100001000111110" => color_data <= "011100110001";
      when "100001000111111" => color_data <= "011100110001";
      when "100001001000000" => color_data <= "011100110001";
      when "100001001000001" => color_data <= "011100110001";
      when "100001001000010" => color_data <= "011100110001";
      when "100001001000011" => color_data <= "011101000001";
      when "100001001000100" => color_data <= "011101000010";
      when "100001001000101" => color_data <= "011000110001";
      when "100001001000110" => color_data <= "011000100000";
      when "100001001000111" => color_data <= "011000100000";
      when "100001001001000" => color_data <= "011000100000";
      when "100001001001001" => color_data <= "010100100000";
      when "100001001001010" => color_data <= "010000010000";
      when "100001001001011" => color_data <= "000000000000";
      when "100001001001100" => color_data <= "000000000000";
      when "100001001001101" => color_data <= "000000000000";
      when "100001001001110" => color_data <= "000000000000";
      when "100001001001111" => color_data <= "000000000000";
      when "100001001010000" => color_data <= "000000000000";
      when "100001001010001" => color_data <= "000000000000";
      when "100001001010010" => color_data <= "000000000000";
      when "100001001010011" => color_data <= "000000000000";
      when "100001001010100" => color_data <= "000000000000";
      when "100001001010101" => color_data <= "000000000000";
      when "100001001010110" => color_data <= "000000000000";
      when "100001001010111" => color_data <= "000000000000";
      when "100001001011000" => color_data <= "000000000000";
      when "100001001011001" => color_data <= "000000000000";
      when "100001001011010" => color_data <= "000000000000";
      when "100001001011011" => color_data <= "000000000000";
      when "100001001011100" => color_data <= "000000000000";
      when "100001001011101" => color_data <= "000000000000";
      when "100001001011110" => color_data <= "000000000000";
      when "100001001011111" => color_data <= "000000000000";
      when "100001001100000" => color_data <= "000000000000";
      when "100001001100001" => color_data <= "000000000000";
      when "100001001100010" => color_data <= "000000000000";
      when "100001001100011" => color_data <= "000000000000";
      when "100001010000000" => color_data <= "000000000000";
      when "100001010000001" => color_data <= "000000000000";
      when "100001010000010" => color_data <= "000000000000";
      when "100001010000011" => color_data <= "000000000000";
      when "100001010000100" => color_data <= "000000000000";
      when "100001010000101" => color_data <= "000000000000";
      when "100001010000110" => color_data <= "000000000000";
      when "100001010000111" => color_data <= "000000000000";
      when "100001010001000" => color_data <= "000000000000";
      when "100001010001001" => color_data <= "000000000000";
      when "100001010001010" => color_data <= "000000000000";
      when "100001010001011" => color_data <= "000000000000";
      when "100001010001100" => color_data <= "000000000000";
      when "100001010001101" => color_data <= "000000000000";
      when "100001010001110" => color_data <= "000000000000";
      when "100001010001111" => color_data <= "000000000000";
      when "100001010010000" => color_data <= "000000000000";
      when "100001010010001" => color_data <= "000000000000";
      when "100001010010010" => color_data <= "000000000000";
      when "100001010010011" => color_data <= "000000000000";
      when "100001010010100" => color_data <= "000000000000";
      when "100001010010101" => color_data <= "000000000000";
      when "100001010010110" => color_data <= "000000000000";
      when "100001010010111" => color_data <= "000000000000";
      when "100001010011000" => color_data <= "000000000000";
      when "100001010011001" => color_data <= "000000000000";
      when "100001010011010" => color_data <= "000000000000";
      when "100001010011011" => color_data <= "010000110011";
      when "100001010011100" => color_data <= "011000100000";
      when "100001010011101" => color_data <= "011101000010";
      when "100001010011110" => color_data <= "011101000001";
      when "100001010011111" => color_data <= "011101000001";
      when "100001010100000" => color_data <= "011101000010";
      when "100001010100001" => color_data <= "011101000001";
      when "100001010100010" => color_data <= "011101000001";
      when "100001010100011" => color_data <= "011101000001";
      when "100001010100100" => color_data <= "011101000001";
      when "100001010100101" => color_data <= "011101000001";
      when "100001010100110" => color_data <= "011101000001";
      when "100001010100111" => color_data <= "011101000001";
      when "100001010101000" => color_data <= "011101000001";
      when "100001010101001" => color_data <= "011101000001";
      when "100001010101010" => color_data <= "011101000001";
      when "100001010101011" => color_data <= "011101000001";
      when "100001010101100" => color_data <= "011101000001";
      when "100001010101101" => color_data <= "011101000001";
      when "100001010101110" => color_data <= "011101000001";
      when "100001010101111" => color_data <= "011101000001";
      when "100001010110000" => color_data <= "011101000001";
      when "100001010110001" => color_data <= "011101000001";
      when "100001010110010" => color_data <= "011101000001";
      when "100001010110011" => color_data <= "011101000001";
      when "100001010110100" => color_data <= "011101000001";
      when "100001010110101" => color_data <= "011101000001";
      when "100001010110110" => color_data <= "011101000001";
      when "100001010110111" => color_data <= "011101000001";
      when "100001010111000" => color_data <= "011101000001";
      when "100001010111001" => color_data <= "011101000001";
      when "100001010111010" => color_data <= "011101000001";
      when "100001010111011" => color_data <= "011101000001";
      when "100001010111100" => color_data <= "011101000001";
      when "100001010111101" => color_data <= "011101000001";
      when "100001010111110" => color_data <= "011101000001";
      when "100001010111111" => color_data <= "011101000001";
      when "100001011000000" => color_data <= "011101000001";
      when "100001011000001" => color_data <= "011101000001";
      when "100001011000010" => color_data <= "011101000001";
      when "100001011000011" => color_data <= "011101000001";
      when "100001011000100" => color_data <= "011101000010";
      when "100001011000101" => color_data <= "011101000010";
      when "100001011000110" => color_data <= "011101000001";
      when "100001011000111" => color_data <= "011101000001";
      when "100001011001000" => color_data <= "011101000001";
      when "100001011001001" => color_data <= "011100110001";
      when "100001011001010" => color_data <= "011000110001";
      when "100001011001011" => color_data <= "000000000000";
      when "100001011001100" => color_data <= "000000000000";
      when "100001011001101" => color_data <= "000000000000";
      when "100001011001110" => color_data <= "000000000000";
      when "100001011001111" => color_data <= "000000000000";
      when "100001011010000" => color_data <= "000000000000";
      when "100001011010001" => color_data <= "000000000000";
      when "100001011010010" => color_data <= "000000000000";
      when "100001011010011" => color_data <= "000000000000";
      when "100001011010100" => color_data <= "000000000000";
      when "100001011010101" => color_data <= "000000000000";
      when "100001011010110" => color_data <= "000000000000";
      when "100001011010111" => color_data <= "000000000000";
      when "100001011011000" => color_data <= "000000000000";
      when "100001011011001" => color_data <= "000000000000";
      when "100001011011010" => color_data <= "000000000000";
      when "100001011011011" => color_data <= "000000000000";
      when "100001011011100" => color_data <= "000000000000";
      when "100001011011101" => color_data <= "000000000000";
      when "100001011011110" => color_data <= "000000000000";
      when "100001011011111" => color_data <= "000000000000";
      when "100001011100000" => color_data <= "000000000000";
      when "100001011100001" => color_data <= "000000000000";
      when "100001011100010" => color_data <= "000000000000";
      when "100001011100011" => color_data <= "000000000000";
      when "100001100000000" => color_data <= "000000000000";
      when "100001100000001" => color_data <= "000000000000";
      when "100001100000010" => color_data <= "000000000000";
      when "100001100000011" => color_data <= "000000000000";
      when "100001100000100" => color_data <= "000000000000";
      when "100001100000101" => color_data <= "000000000000";
      when "100001100000110" => color_data <= "000000000000";
      when "100001100000111" => color_data <= "000000000000";
      when "100001100001000" => color_data <= "000000000000";
      when "100001100001001" => color_data <= "000000000000";
      when "100001100001010" => color_data <= "000000000000";
      when "100001100001011" => color_data <= "000000000000";
      when "100001100001100" => color_data <= "000000000000";
      when "100001100001101" => color_data <= "000000000000";
      when "100001100001110" => color_data <= "000000000000";
      when "100001100001111" => color_data <= "000000000000";
      when "100001100010000" => color_data <= "000000000000";
      when "100001100010001" => color_data <= "000000000000";
      when "100001100010010" => color_data <= "000000000000";
      when "100001100010011" => color_data <= "000000000000";
      when "100001100010100" => color_data <= "000000000000";
      when "100001100010101" => color_data <= "000000000000";
      when "100001100010110" => color_data <= "000000000000";
      when "100001100010111" => color_data <= "000000000000";
      when "100001100011000" => color_data <= "000000000000";
      when "100001100011001" => color_data <= "000000000000";
      when "100001100011010" => color_data <= "000000000000";
      when "100001100011011" => color_data <= "010000110011";
      when "100001100011100" => color_data <= "011000100000";
      when "100001100011101" => color_data <= "011101000010";
      when "100001100011110" => color_data <= "011101000010";
      when "100001100011111" => color_data <= "011101000001";
      when "100001100100000" => color_data <= "011000100000";
      when "100001100100001" => color_data <= "101010000101";
      when "100001100100010" => color_data <= "111011101001";
      when "100001100100011" => color_data <= "111011001000";
      when "100001100100100" => color_data <= "111011001000";
      when "100001100100101" => color_data <= "111011001000";
      when "100001100100110" => color_data <= "111011001000";
      when "100001100100111" => color_data <= "111011001000";
      when "100001100101000" => color_data <= "111011001000";
      when "100001100101001" => color_data <= "111011001000";
      when "100001100101010" => color_data <= "111011001000";
      when "100001100101011" => color_data <= "111011001000";
      when "100001100101100" => color_data <= "111011001000";
      when "100001100101101" => color_data <= "111011001000";
      when "100001100101110" => color_data <= "111011001000";
      when "100001100101111" => color_data <= "111011001000";
      when "100001100110000" => color_data <= "111011001000";
      when "100001100110001" => color_data <= "111011001000";
      when "100001100110010" => color_data <= "111011001000";
      when "100001100110011" => color_data <= "111011001000";
      when "100001100110100" => color_data <= "111011001000";
      when "100001100110101" => color_data <= "111011001000";
      when "100001100110110" => color_data <= "111011001000";
      when "100001100110111" => color_data <= "111011001000";
      when "100001100111000" => color_data <= "111011001000";
      when "100001100111001" => color_data <= "111011001000";
      when "100001100111010" => color_data <= "111011001000";
      when "100001100111011" => color_data <= "111011001000";
      when "100001100111100" => color_data <= "111011001000";
      when "100001100111101" => color_data <= "111011001000";
      when "100001100111110" => color_data <= "111011001000";
      when "100001100111111" => color_data <= "111011001000";
      when "100001101000000" => color_data <= "111011001000";
      when "100001101000001" => color_data <= "111011001000";
      when "100001101000010" => color_data <= "111011101001";
      when "100001101000011" => color_data <= "101110100110";
      when "100001101000100" => color_data <= "011000110001";
      when "100001101000101" => color_data <= "011101000010";
      when "100001101000110" => color_data <= "011101000010";
      when "100001101000111" => color_data <= "011101000010";
      when "100001101001000" => color_data <= "011101000010";
      when "100001101001001" => color_data <= "011100110001";
      when "100001101001010" => color_data <= "011000110001";
      when "100001101001011" => color_data <= "000000000000";
      when "100001101001100" => color_data <= "000000000000";
      when "100001101001101" => color_data <= "000000000000";
      when "100001101001110" => color_data <= "000000000000";
      when "100001101001111" => color_data <= "000000000000";
      when "100001101010000" => color_data <= "000000000000";
      when "100001101010001" => color_data <= "000000000000";
      when "100001101010010" => color_data <= "000000000000";
      when "100001101010011" => color_data <= "000000000000";
      when "100001101010100" => color_data <= "000000000000";
      when "100001101010101" => color_data <= "000000000000";
      when "100001101010110" => color_data <= "000000000000";
      when "100001101010111" => color_data <= "000000000000";
      when "100001101011000" => color_data <= "000000000000";
      when "100001101011001" => color_data <= "000000000000";
      when "100001101011010" => color_data <= "000000000000";
      when "100001101011011" => color_data <= "000000000000";
      when "100001101011100" => color_data <= "000000000000";
      when "100001101011101" => color_data <= "000000000000";
      when "100001101011110" => color_data <= "000000000000";
      when "100001101011111" => color_data <= "000000000000";
      when "100001101100000" => color_data <= "000000000000";
      when "100001101100001" => color_data <= "000000000000";
      when "100001101100010" => color_data <= "000000000000";
      when "100001101100011" => color_data <= "000000000000";
      when "100001110000000" => color_data <= "000000000000";
      when "100001110000001" => color_data <= "000000000000";
      when "100001110000010" => color_data <= "000000000000";
      when "100001110000011" => color_data <= "000000000000";
      when "100001110000100" => color_data <= "000000000000";
      when "100001110000101" => color_data <= "000000000000";
      when "100001110000110" => color_data <= "000000000000";
      when "100001110000111" => color_data <= "000000000000";
      when "100001110001000" => color_data <= "000000000000";
      when "100001110001001" => color_data <= "000000000000";
      when "100001110001010" => color_data <= "000000000000";
      when "100001110001011" => color_data <= "000000000000";
      when "100001110001100" => color_data <= "000000000000";
      when "100001110001101" => color_data <= "000000000000";
      when "100001110001110" => color_data <= "000000000000";
      when "100001110001111" => color_data <= "000000000000";
      when "100001110010000" => color_data <= "000000000000";
      when "100001110010001" => color_data <= "000000000000";
      when "100001110010010" => color_data <= "000000000000";
      when "100001110010011" => color_data <= "000000000000";
      when "100001110010100" => color_data <= "000000000000";
      when "100001110010101" => color_data <= "000000000000";
      when "100001110010110" => color_data <= "000000000000";
      when "100001110010111" => color_data <= "000000000000";
      when "100001110011000" => color_data <= "000000000000";
      when "100001110011001" => color_data <= "000000000000";
      when "100001110011010" => color_data <= "000000000000";
      when "100001110011011" => color_data <= "010000110011";
      when "100001110011100" => color_data <= "011000100000";
      when "100001110011101" => color_data <= "011101000010";
      when "100001110011110" => color_data <= "011101000010";
      when "100001110011111" => color_data <= "011101000010";
      when "100001110100000" => color_data <= "010100100000";
      when "100001110100001" => color_data <= "101110010101";
      when "100001110100010" => color_data <= "111111111100";
      when "100001110100011" => color_data <= "111111111010";
      when "100001110100100" => color_data <= "111111111010";
      when "100001110100101" => color_data <= "111111111010";
      when "100001110100110" => color_data <= "111111111010";
      when "100001110100111" => color_data <= "111111111010";
      when "100001110101000" => color_data <= "111111111010";
      when "100001110101001" => color_data <= "111111111010";
      when "100001110101010" => color_data <= "111111111010";
      when "100001110101011" => color_data <= "111111111010";
      when "100001110101100" => color_data <= "111111111010";
      when "100001110101101" => color_data <= "111111111010";
      when "100001110101110" => color_data <= "111111111010";
      when "100001110101111" => color_data <= "111111111010";
      when "100001110110000" => color_data <= "111111111010";
      when "100001110110001" => color_data <= "111111111010";
      when "100001110110010" => color_data <= "111111111010";
      when "100001110110011" => color_data <= "111111111010";
      when "100001110110100" => color_data <= "111111111010";
      when "100001110110101" => color_data <= "111111111010";
      when "100001110110110" => color_data <= "111111111010";
      when "100001110110111" => color_data <= "111111111010";
      when "100001110111000" => color_data <= "111111111010";
      when "100001110111001" => color_data <= "111111111010";
      when "100001110111010" => color_data <= "111111111010";
      when "100001110111011" => color_data <= "111111111010";
      when "100001110111100" => color_data <= "111111111010";
      when "100001110111101" => color_data <= "111111111010";
      when "100001110111110" => color_data <= "111111111010";
      when "100001110111111" => color_data <= "111111111010";
      when "100001111000000" => color_data <= "111111111010";
      when "100001111000001" => color_data <= "111111111010";
      when "100001111000010" => color_data <= "111111111011";
      when "100001111000011" => color_data <= "110110110111";
      when "100001111000100" => color_data <= "011000100000";
      when "100001111000101" => color_data <= "011101000010";
      when "100001111000110" => color_data <= "011101000010";
      when "100001111000111" => color_data <= "011101000010";
      when "100001111001000" => color_data <= "011101000010";
      when "100001111001001" => color_data <= "011100110001";
      when "100001111001010" => color_data <= "011000110001";
      when "100001111001011" => color_data <= "000000000000";
      when "100001111001100" => color_data <= "000000000000";
      when "100001111001101" => color_data <= "000000000000";
      when "100001111001110" => color_data <= "000000000000";
      when "100001111001111" => color_data <= "000000000000";
      when "100001111010000" => color_data <= "000000000000";
      when "100001111010001" => color_data <= "000000000000";
      when "100001111010010" => color_data <= "000000000000";
      when "100001111010011" => color_data <= "000000000000";
      when "100001111010100" => color_data <= "000000000000";
      when "100001111010101" => color_data <= "000000000000";
      when "100001111010110" => color_data <= "000000000000";
      when "100001111010111" => color_data <= "000000000000";
      when "100001111011000" => color_data <= "000000000000";
      when "100001111011001" => color_data <= "000000000000";
      when "100001111011010" => color_data <= "000000000000";
      when "100001111011011" => color_data <= "000000000000";
      when "100001111011100" => color_data <= "000000000000";
      when "100001111011101" => color_data <= "000000000000";
      when "100001111011110" => color_data <= "000000000000";
      when "100001111011111" => color_data <= "000000000000";
      when "100001111100000" => color_data <= "000000000000";
      when "100001111100001" => color_data <= "000000000000";
      when "100001111100010" => color_data <= "000000000000";
      when "100001111100011" => color_data <= "000000000000";
      when "100010000000000" => color_data <= "000000000000";
      when "100010000000001" => color_data <= "000000000000";
      when "100010000000010" => color_data <= "000000000000";
      when "100010000000011" => color_data <= "000000000000";
      when "100010000000100" => color_data <= "000000000000";
      when "100010000000101" => color_data <= "000000000000";
      when "100010000000110" => color_data <= "000000000000";
      when "100010000000111" => color_data <= "000000000000";
      when "100010000001000" => color_data <= "000000000000";
      when "100010000001001" => color_data <= "000000000000";
      when "100010000001010" => color_data <= "000000000000";
      when "100010000001011" => color_data <= "000000000000";
      when "100010000001100" => color_data <= "000000000000";
      when "100010000001101" => color_data <= "000000000000";
      when "100010000001110" => color_data <= "000000000000";
      when "100010000001111" => color_data <= "000000000000";
      when "100010000010000" => color_data <= "000000000000";
      when "100010000010001" => color_data <= "000000000000";
      when "100010000010010" => color_data <= "000000000000";
      when "100010000010011" => color_data <= "000000000000";
      when "100010000010100" => color_data <= "000000000000";
      when "100010000010101" => color_data <= "000000000000";
      when "100010000010110" => color_data <= "000000000000";
      when "100010000010111" => color_data <= "000000000000";
      when "100010000011000" => color_data <= "000000000000";
      when "100010000011001" => color_data <= "000000000000";
      when "100010000011010" => color_data <= "000000000000";
      when "100010000011011" => color_data <= "010000110011";
      when "100010000011100" => color_data <= "011000100000";
      when "100010000011101" => color_data <= "011101000010";
      when "100010000011110" => color_data <= "011101000010";
      when "100010000011111" => color_data <= "011101000010";
      when "100010000100000" => color_data <= "011000100000";
      when "100010000100001" => color_data <= "101110010101";
      when "100010000100010" => color_data <= "111111111011";
      when "100010000100011" => color_data <= "111111101001";
      when "100010000100100" => color_data <= "111111101001";
      when "100010000100101" => color_data <= "111111101001";
      when "100010000100110" => color_data <= "111111101001";
      when "100010000100111" => color_data <= "111111101001";
      when "100010000101000" => color_data <= "111111101001";
      when "100010000101001" => color_data <= "111111101001";
      when "100010000101010" => color_data <= "111111101001";
      when "100010000101011" => color_data <= "111111101001";
      when "100010000101100" => color_data <= "111111101001";
      when "100010000101101" => color_data <= "111111101001";
      when "100010000101110" => color_data <= "111111101001";
      when "100010000101111" => color_data <= "111111101001";
      when "100010000110000" => color_data <= "111111101001";
      when "100010000110001" => color_data <= "111111101001";
      when "100010000110010" => color_data <= "111111101001";
      when "100010000110011" => color_data <= "111111101001";
      when "100010000110100" => color_data <= "111111101001";
      when "100010000110101" => color_data <= "111111101001";
      when "100010000110110" => color_data <= "111111101001";
      when "100010000110111" => color_data <= "111111101001";
      when "100010000111000" => color_data <= "111111101001";
      when "100010000111001" => color_data <= "111111101001";
      when "100010000111010" => color_data <= "111111101001";
      when "100010000111011" => color_data <= "111111101001";
      when "100010000111100" => color_data <= "111111101001";
      when "100010000111101" => color_data <= "111111101001";
      when "100010000111110" => color_data <= "111111101001";
      when "100010000111111" => color_data <= "111111101001";
      when "100010001000000" => color_data <= "111111101001";
      when "100010001000001" => color_data <= "111111101001";
      when "100010001000010" => color_data <= "111111111010";
      when "100010001000011" => color_data <= "110010110110";
      when "100010001000100" => color_data <= "011000100000";
      when "100010001000101" => color_data <= "011101000010";
      when "100010001000110" => color_data <= "011101000010";
      when "100010001000111" => color_data <= "011101000010";
      when "100010001001000" => color_data <= "011101000010";
      when "100010001001001" => color_data <= "011100110001";
      when "100010001001010" => color_data <= "011000110001";
      when "100010001001011" => color_data <= "000000000000";
      when "100010001001100" => color_data <= "000000000000";
      when "100010001001101" => color_data <= "000000000000";
      when "100010001001110" => color_data <= "000000000000";
      when "100010001001111" => color_data <= "000000000000";
      when "100010001010000" => color_data <= "000000000000";
      when "100010001010001" => color_data <= "000000000000";
      when "100010001010010" => color_data <= "000000000000";
      when "100010001010011" => color_data <= "000000000000";
      when "100010001010100" => color_data <= "000000000000";
      when "100010001010101" => color_data <= "000000000000";
      when "100010001010110" => color_data <= "000000000000";
      when "100010001010111" => color_data <= "000000000000";
      when "100010001011000" => color_data <= "000000000000";
      when "100010001011001" => color_data <= "000000000000";
      when "100010001011010" => color_data <= "000000000000";
      when "100010001011011" => color_data <= "000000000000";
      when "100010001011100" => color_data <= "000000000000";
      when "100010001011101" => color_data <= "000000000000";
      when "100010001011110" => color_data <= "000000000000";
      when "100010001011111" => color_data <= "000000000000";
      when "100010001100000" => color_data <= "000000000000";
      when "100010001100001" => color_data <= "000000000000";
      when "100010001100010" => color_data <= "000000000000";
      when "100010001100011" => color_data <= "000000000000";
      when "100010010000000" => color_data <= "000000000000";
      when "100010010000001" => color_data <= "000000000000";
      when "100010010000010" => color_data <= "000000000000";
      when "100010010000011" => color_data <= "000000000000";
      when "100010010000100" => color_data <= "000000000000";
      when "100010010000101" => color_data <= "000000000000";
      when "100010010000110" => color_data <= "000000000000";
      when "100010010000111" => color_data <= "000000000000";
      when "100010010001000" => color_data <= "000000000000";
      when "100010010001001" => color_data <= "000000000000";
      when "100010010001010" => color_data <= "000000000000";
      when "100010010001011" => color_data <= "000000000000";
      when "100010010001100" => color_data <= "000000000000";
      when "100010010001101" => color_data <= "000000000000";
      when "100010010001110" => color_data <= "000000000000";
      when "100010010001111" => color_data <= "000000000000";
      when "100010010010000" => color_data <= "000000000000";
      when "100010010010001" => color_data <= "000000000000";
      when "100010010010010" => color_data <= "000000000000";
      when "100010010010011" => color_data <= "000000000000";
      when "100010010010100" => color_data <= "000000000000";
      when "100010010010101" => color_data <= "000000000000";
      when "100010010010110" => color_data <= "000000000000";
      when "100010010010111" => color_data <= "000000000000";
      when "100010010011000" => color_data <= "000000000000";
      when "100010010011001" => color_data <= "000000000000";
      when "100010010011010" => color_data <= "000000000000";
      when "100010010011011" => color_data <= "010000110011";
      when "100010010011100" => color_data <= "011000100000";
      when "100010010011101" => color_data <= "011101000010";
      when "100010010011110" => color_data <= "011101000010";
      when "100010010011111" => color_data <= "011101000010";
      when "100010010100000" => color_data <= "011000100000";
      when "100010010100001" => color_data <= "101110010101";
      when "100010010100010" => color_data <= "111111111011";
      when "100010010100011" => color_data <= "111111101001";
      when "100010010100100" => color_data <= "111111101001";
      when "100010010100101" => color_data <= "111111101001";
      when "100010010100110" => color_data <= "111111101001";
      when "100010010100111" => color_data <= "111111101001";
      when "100010010101000" => color_data <= "111111101001";
      when "100010010101001" => color_data <= "111111101001";
      when "100010010101010" => color_data <= "111111101001";
      when "100010010101011" => color_data <= "111111101001";
      when "100010010101100" => color_data <= "111111101001";
      when "100010010101101" => color_data <= "111111101001";
      when "100010010101110" => color_data <= "111111101001";
      when "100010010101111" => color_data <= "111111101001";
      when "100010010110000" => color_data <= "111111101001";
      when "100010010110001" => color_data <= "111111101001";
      when "100010010110010" => color_data <= "111111101001";
      when "100010010110011" => color_data <= "111111101001";
      when "100010010110100" => color_data <= "111111101001";
      when "100010010110101" => color_data <= "111111101001";
      when "100010010110110" => color_data <= "111111101001";
      when "100010010110111" => color_data <= "111111101001";
      when "100010010111000" => color_data <= "111111101001";
      when "100010010111001" => color_data <= "111111101001";
      when "100010010111010" => color_data <= "111111101001";
      when "100010010111011" => color_data <= "111111101001";
      when "100010010111100" => color_data <= "111111101001";
      when "100010010111101" => color_data <= "111111101001";
      when "100010010111110" => color_data <= "111111101001";
      when "100010010111111" => color_data <= "111111101001";
      when "100010011000000" => color_data <= "111111101001";
      when "100010011000001" => color_data <= "111111101001";
      when "100010011000010" => color_data <= "111111111010";
      when "100010011000011" => color_data <= "110010110110";
      when "100010011000100" => color_data <= "011000100000";
      when "100010011000101" => color_data <= "011101000010";
      when "100010011000110" => color_data <= "011101000010";
      when "100010011000111" => color_data <= "011101000010";
      when "100010011001000" => color_data <= "011101000010";
      when "100010011001001" => color_data <= "011100110001";
      when "100010011001010" => color_data <= "011000110001";
      when "100010011001011" => color_data <= "000000000000";
      when "100010011001100" => color_data <= "000000000000";
      when "100010011001101" => color_data <= "000000000000";
      when "100010011001110" => color_data <= "000000000000";
      when "100010011001111" => color_data <= "000000000000";
      when "100010011010000" => color_data <= "000000000000";
      when "100010011010001" => color_data <= "000000000000";
      when "100010011010010" => color_data <= "000000000000";
      when "100010011010011" => color_data <= "000000000000";
      when "100010011010100" => color_data <= "000000000000";
      when "100010011010101" => color_data <= "000000000000";
      when "100010011010110" => color_data <= "000000000000";
      when "100010011010111" => color_data <= "000000000000";
      when "100010011011000" => color_data <= "000000000000";
      when "100010011011001" => color_data <= "000000000000";
      when "100010011011010" => color_data <= "000000000000";
      when "100010011011011" => color_data <= "000000000000";
      when "100010011011100" => color_data <= "000000000000";
      when "100010011011101" => color_data <= "000000000000";
      when "100010011011110" => color_data <= "000000000000";
      when "100010011011111" => color_data <= "000000000000";
      when "100010011100000" => color_data <= "000000000000";
      when "100010011100001" => color_data <= "000000000000";
      when "100010011100010" => color_data <= "000000000000";
      when "100010011100011" => color_data <= "000000000000";
      when "100010100000000" => color_data <= "000000000000";
      when "100010100000001" => color_data <= "000000000000";
      when "100010100000010" => color_data <= "000000000000";
      when "100010100000011" => color_data <= "000000000000";
      when "100010100000100" => color_data <= "000000000000";
      when "100010100000101" => color_data <= "000000000000";
      when "100010100000110" => color_data <= "000000000000";
      when "100010100000111" => color_data <= "000000000000";
      when "100010100001000" => color_data <= "000000000000";
      when "100010100001001" => color_data <= "000000000000";
      when "100010100001010" => color_data <= "000000000000";
      when "100010100001011" => color_data <= "000000000000";
      when "100010100001100" => color_data <= "000000000000";
      when "100010100001101" => color_data <= "000000000000";
      when "100010100001110" => color_data <= "000000000000";
      when "100010100001111" => color_data <= "000000000000";
      when "100010100010000" => color_data <= "000000000000";
      when "100010100010001" => color_data <= "000000000000";
      when "100010100010010" => color_data <= "000000000000";
      when "100010100010011" => color_data <= "000000000000";
      when "100010100010100" => color_data <= "000000000000";
      when "100010100010101" => color_data <= "000000000000";
      when "100010100010110" => color_data <= "000000000000";
      when "100010100010111" => color_data <= "000000000000";
      when "100010100011000" => color_data <= "000000000000";
      when "100010100011001" => color_data <= "000000000000";
      when "100010100011010" => color_data <= "000000000000";
      when "100010100011011" => color_data <= "010000110011";
      when "100010100011100" => color_data <= "011000100000";
      when "100010100011101" => color_data <= "011101000010";
      when "100010100011110" => color_data <= "011101000010";
      when "100010100011111" => color_data <= "011101000010";
      when "100010100100000" => color_data <= "011000100000";
      when "100010100100001" => color_data <= "101110010101";
      when "100010100100010" => color_data <= "111111111011";
      when "100010100100011" => color_data <= "111111101001";
      when "100010100100100" => color_data <= "111111101001";
      when "100010100100101" => color_data <= "111111101001";
      when "100010100100110" => color_data <= "111111101001";
      when "100010100100111" => color_data <= "111111101001";
      when "100010100101000" => color_data <= "111111101001";
      when "100010100101001" => color_data <= "111111101001";
      when "100010100101010" => color_data <= "111111101001";
      when "100010100101011" => color_data <= "111111101001";
      when "100010100101100" => color_data <= "111111101001";
      when "100010100101101" => color_data <= "111111101001";
      when "100010100101110" => color_data <= "111111101001";
      when "100010100101111" => color_data <= "111111101001";
      when "100010100110000" => color_data <= "111111101001";
      when "100010100110001" => color_data <= "111111101001";
      when "100010100110010" => color_data <= "111111101001";
      when "100010100110011" => color_data <= "111111101001";
      when "100010100110100" => color_data <= "111111101001";
      when "100010100110101" => color_data <= "111111101001";
      when "100010100110110" => color_data <= "111111101001";
      when "100010100110111" => color_data <= "111111101001";
      when "100010100111000" => color_data <= "111111101001";
      when "100010100111001" => color_data <= "111111101001";
      when "100010100111010" => color_data <= "111111101001";
      when "100010100111011" => color_data <= "111111101001";
      when "100010100111100" => color_data <= "111111101001";
      when "100010100111101" => color_data <= "111111101001";
      when "100010100111110" => color_data <= "111111101001";
      when "100010100111111" => color_data <= "111111101001";
      when "100010101000000" => color_data <= "111111101001";
      when "100010101000001" => color_data <= "111111101001";
      when "100010101000010" => color_data <= "111111111010";
      when "100010101000011" => color_data <= "110010110110";
      when "100010101000100" => color_data <= "011000100000";
      when "100010101000101" => color_data <= "011101000010";
      when "100010101000110" => color_data <= "011101000010";
      when "100010101000111" => color_data <= "011101000010";
      when "100010101001000" => color_data <= "011101000010";
      when "100010101001001" => color_data <= "011100110001";
      when "100010101001010" => color_data <= "011000110001";
      when "100010101001011" => color_data <= "000000000000";
      when "100010101001100" => color_data <= "000000000000";
      when "100010101001101" => color_data <= "000000000000";
      when "100010101001110" => color_data <= "000000000000";
      when "100010101001111" => color_data <= "000000000000";
      when "100010101010000" => color_data <= "000000000000";
      when "100010101010001" => color_data <= "000000000000";
      when "100010101010010" => color_data <= "000000000000";
      when "100010101010011" => color_data <= "000000000000";
      when "100010101010100" => color_data <= "000000000000";
      when "100010101010101" => color_data <= "000000000000";
      when "100010101010110" => color_data <= "000000000000";
      when "100010101010111" => color_data <= "000000000000";
      when "100010101011000" => color_data <= "000000000000";
      when "100010101011001" => color_data <= "000000000000";
      when "100010101011010" => color_data <= "000000000000";
      when "100010101011011" => color_data <= "000000000000";
      when "100010101011100" => color_data <= "000000000000";
      when "100010101011101" => color_data <= "000000000000";
      when "100010101011110" => color_data <= "000000000000";
      when "100010101011111" => color_data <= "000000000000";
      when "100010101100000" => color_data <= "000000000000";
      when "100010101100001" => color_data <= "000000000000";
      when "100010101100010" => color_data <= "000000000000";
      when "100010101100011" => color_data <= "000000000000";
      when "100010110000000" => color_data <= "000000000000";
      when "100010110000001" => color_data <= "000000000000";
      when "100010110000010" => color_data <= "000000000000";
      when "100010110000011" => color_data <= "000000000000";
      when "100010110000100" => color_data <= "000000000000";
      when "100010110000101" => color_data <= "000000000000";
      when "100010110000110" => color_data <= "000000000000";
      when "100010110000111" => color_data <= "000000000000";
      when "100010110001000" => color_data <= "000000000000";
      when "100010110001001" => color_data <= "000000000000";
      when "100010110001010" => color_data <= "000000000000";
      when "100010110001011" => color_data <= "000000000000";
      when "100010110001100" => color_data <= "000000000000";
      when "100010110001101" => color_data <= "000000000000";
      when "100010110001110" => color_data <= "000000000000";
      when "100010110001111" => color_data <= "000000000000";
      when "100010110010000" => color_data <= "000000000000";
      when "100010110010001" => color_data <= "000000000000";
      when "100010110010010" => color_data <= "000000000000";
      when "100010110010011" => color_data <= "000000000000";
      when "100010110010100" => color_data <= "000000000000";
      when "100010110010101" => color_data <= "000000000000";
      when "100010110010110" => color_data <= "000000000000";
      when "100010110010111" => color_data <= "000000000000";
      when "100010110011000" => color_data <= "000000000000";
      when "100010110011001" => color_data <= "000000000000";
      when "100010110011010" => color_data <= "000000000000";
      when "100010110011011" => color_data <= "010000110011";
      when "100010110011100" => color_data <= "011000100000";
      when "100010110011101" => color_data <= "011101000010";
      when "100010110011110" => color_data <= "011101000010";
      when "100010110011111" => color_data <= "011101000010";
      when "100010110100000" => color_data <= "011000100000";
      when "100010110100001" => color_data <= "101110010101";
      when "100010110100010" => color_data <= "111111111011";
      when "100010110100011" => color_data <= "111111101001";
      when "100010110100100" => color_data <= "111111101001";
      when "100010110100101" => color_data <= "111111101001";
      when "100010110100110" => color_data <= "111111101001";
      when "100010110100111" => color_data <= "111111101001";
      when "100010110101000" => color_data <= "111111101001";
      when "100010110101001" => color_data <= "111111101001";
      when "100010110101010" => color_data <= "111111101001";
      when "100010110101011" => color_data <= "111111101001";
      when "100010110101100" => color_data <= "111111101001";
      when "100010110101101" => color_data <= "111111101001";
      when "100010110101110" => color_data <= "111111101001";
      when "100010110101111" => color_data <= "111111101001";
      when "100010110110000" => color_data <= "111111101001";
      when "100010110110001" => color_data <= "111111101001";
      when "100010110110010" => color_data <= "111111101001";
      when "100010110110011" => color_data <= "111111101001";
      when "100010110110100" => color_data <= "111111101001";
      when "100010110110101" => color_data <= "111111101001";
      when "100010110110110" => color_data <= "111111101001";
      when "100010110110111" => color_data <= "111111101001";
      when "100010110111000" => color_data <= "111111101001";
      when "100010110111001" => color_data <= "111111101001";
      when "100010110111010" => color_data <= "111111101001";
      when "100010110111011" => color_data <= "111111101001";
      when "100010110111100" => color_data <= "111111101001";
      when "100010110111101" => color_data <= "111111101001";
      when "100010110111110" => color_data <= "111111101001";
      when "100010110111111" => color_data <= "111111101001";
      when "100010111000000" => color_data <= "111111101001";
      when "100010111000001" => color_data <= "111111101001";
      when "100010111000010" => color_data <= "111111111010";
      when "100010111000011" => color_data <= "110010110110";
      when "100010111000100" => color_data <= "011000100000";
      when "100010111000101" => color_data <= "011101000010";
      when "100010111000110" => color_data <= "011101000010";
      when "100010111000111" => color_data <= "011101000010";
      when "100010111001000" => color_data <= "011101000010";
      when "100010111001001" => color_data <= "011100110001";
      when "100010111001010" => color_data <= "011000110001";
      when "100010111001011" => color_data <= "000000000000";
      when "100010111001100" => color_data <= "000000000000";
      when "100010111001101" => color_data <= "000000000000";
      when "100010111001110" => color_data <= "000000000000";
      when "100010111001111" => color_data <= "000000000000";
      when "100010111010000" => color_data <= "000000000000";
      when "100010111010001" => color_data <= "000000000000";
      when "100010111010010" => color_data <= "000000000000";
      when "100010111010011" => color_data <= "000000000000";
      when "100010111010100" => color_data <= "000000000000";
      when "100010111010101" => color_data <= "000000000000";
      when "100010111010110" => color_data <= "000000000000";
      when "100010111010111" => color_data <= "000000000000";
      when "100010111011000" => color_data <= "000000000000";
      when "100010111011001" => color_data <= "000000000000";
      when "100010111011010" => color_data <= "000000000000";
      when "100010111011011" => color_data <= "000000000000";
      when "100010111011100" => color_data <= "000000000000";
      when "100010111011101" => color_data <= "000000000000";
      when "100010111011110" => color_data <= "000000000000";
      when "100010111011111" => color_data <= "000000000000";
      when "100010111100000" => color_data <= "000000000000";
      when "100010111100001" => color_data <= "000000000000";
      when "100010111100010" => color_data <= "000000000000";
      when "100010111100011" => color_data <= "000000000000";
      when "100011000000000" => color_data <= "000000000000";
      when "100011000000001" => color_data <= "000000000000";
      when "100011000000010" => color_data <= "000000000000";
      when "100011000000011" => color_data <= "000000000000";
      when "100011000000100" => color_data <= "000000000000";
      when "100011000000101" => color_data <= "000000000000";
      when "100011000000110" => color_data <= "000000000000";
      when "100011000000111" => color_data <= "000000000000";
      when "100011000001000" => color_data <= "000000000000";
      when "100011000001001" => color_data <= "000000000000";
      when "100011000001010" => color_data <= "000000000000";
      when "100011000001011" => color_data <= "000000000000";
      when "100011000001100" => color_data <= "000000000000";
      when "100011000001101" => color_data <= "000000000000";
      when "100011000001110" => color_data <= "000000000000";
      when "100011000001111" => color_data <= "000000000000";
      when "100011000010000" => color_data <= "000000000000";
      when "100011000010001" => color_data <= "000000000000";
      when "100011000010010" => color_data <= "000000000000";
      when "100011000010011" => color_data <= "000000000000";
      when "100011000010100" => color_data <= "000000000000";
      when "100011000010101" => color_data <= "000000000000";
      when "100011000010110" => color_data <= "000000000000";
      when "100011000010111" => color_data <= "000000000000";
      when "100011000011000" => color_data <= "000000000000";
      when "100011000011001" => color_data <= "000000000000";
      when "100011000011010" => color_data <= "000000000000";
      when "100011000011011" => color_data <= "010000110011";
      when "100011000011100" => color_data <= "011000100000";
      when "100011000011101" => color_data <= "011101000010";
      when "100011000011110" => color_data <= "011101000010";
      when "100011000011111" => color_data <= "011101000010";
      when "100011000100000" => color_data <= "011000100000";
      when "100011000100001" => color_data <= "101110010101";
      when "100011000100010" => color_data <= "111111111011";
      when "100011000100011" => color_data <= "111111101001";
      when "100011000100100" => color_data <= "111111101001";
      when "100011000100101" => color_data <= "111111101001";
      when "100011000100110" => color_data <= "111111101001";
      when "100011000100111" => color_data <= "111111101001";
      when "100011000101000" => color_data <= "111111101001";
      when "100011000101001" => color_data <= "111111101001";
      when "100011000101010" => color_data <= "111111101001";
      when "100011000101011" => color_data <= "111111101001";
      when "100011000101100" => color_data <= "111111101001";
      when "100011000101101" => color_data <= "111111101001";
      when "100011000101110" => color_data <= "111111101001";
      when "100011000101111" => color_data <= "111111101001";
      when "100011000110000" => color_data <= "111111101001";
      when "100011000110001" => color_data <= "111111101001";
      when "100011000110010" => color_data <= "111111101001";
      when "100011000110011" => color_data <= "111111101001";
      when "100011000110100" => color_data <= "111111101001";
      when "100011000110101" => color_data <= "111111101001";
      when "100011000110110" => color_data <= "111111101001";
      when "100011000110111" => color_data <= "111111101001";
      when "100011000111000" => color_data <= "111111101001";
      when "100011000111001" => color_data <= "111111101001";
      when "100011000111010" => color_data <= "111111101001";
      when "100011000111011" => color_data <= "111111101001";
      when "100011000111100" => color_data <= "111111101001";
      when "100011000111101" => color_data <= "111111101001";
      when "100011000111110" => color_data <= "111111101001";
      when "100011000111111" => color_data <= "111111101001";
      when "100011001000000" => color_data <= "111111101001";
      when "100011001000001" => color_data <= "111111101001";
      when "100011001000010" => color_data <= "111111111010";
      when "100011001000011" => color_data <= "110010110110";
      when "100011001000100" => color_data <= "011000100000";
      when "100011001000101" => color_data <= "011101000010";
      when "100011001000110" => color_data <= "011101000010";
      when "100011001000111" => color_data <= "011101000010";
      when "100011001001000" => color_data <= "011101000010";
      when "100011001001001" => color_data <= "011100110001";
      when "100011001001010" => color_data <= "011000110001";
      when "100011001001011" => color_data <= "000000000000";
      when "100011001001100" => color_data <= "000000000000";
      when "100011001001101" => color_data <= "000000000000";
      when "100011001001110" => color_data <= "000000000000";
      when "100011001001111" => color_data <= "000000000000";
      when "100011001010000" => color_data <= "000000000000";
      when "100011001010001" => color_data <= "000000000000";
      when "100011001010010" => color_data <= "000000000000";
      when "100011001010011" => color_data <= "000000000000";
      when "100011001010100" => color_data <= "000000000000";
      when "100011001010101" => color_data <= "000000000000";
      when "100011001010110" => color_data <= "000000000000";
      when "100011001010111" => color_data <= "000000000000";
      when "100011001011000" => color_data <= "000000000000";
      when "100011001011001" => color_data <= "000000000000";
      when "100011001011010" => color_data <= "000000000000";
      when "100011001011011" => color_data <= "000000000000";
      when "100011001011100" => color_data <= "000000000000";
      when "100011001011101" => color_data <= "000000000000";
      when "100011001011110" => color_data <= "000000000000";
      when "100011001011111" => color_data <= "000000000000";
      when "100011001100000" => color_data <= "000000000000";
      when "100011001100001" => color_data <= "000000000000";
      when "100011001100010" => color_data <= "000000000000";
      when "100011001100011" => color_data <= "000000000000";
      when "100011010000000" => color_data <= "000000000000";
      when "100011010000001" => color_data <= "000000000000";
      when "100011010000010" => color_data <= "000000000000";
      when "100011010000011" => color_data <= "000000000000";
      when "100011010000100" => color_data <= "000000000000";
      when "100011010000101" => color_data <= "000000000000";
      when "100011010000110" => color_data <= "000000000000";
      when "100011010000111" => color_data <= "000000000000";
      when "100011010001000" => color_data <= "000000000000";
      when "100011010001001" => color_data <= "000000000000";
      when "100011010001010" => color_data <= "000000000000";
      when "100011010001011" => color_data <= "000000000000";
      when "100011010001100" => color_data <= "000000000000";
      when "100011010001101" => color_data <= "000000000000";
      when "100011010001110" => color_data <= "000000000000";
      when "100011010001111" => color_data <= "000000000000";
      when "100011010010000" => color_data <= "000000000000";
      when "100011010010001" => color_data <= "000000000000";
      when "100011010010010" => color_data <= "000000000000";
      when "100011010010011" => color_data <= "000000000000";
      when "100011010010100" => color_data <= "000000000000";
      when "100011010010101" => color_data <= "000000000000";
      when "100011010010110" => color_data <= "000000000000";
      when "100011010010111" => color_data <= "000000000000";
      when "100011010011000" => color_data <= "000000000000";
      when "100011010011001" => color_data <= "000000000000";
      when "100011010011010" => color_data <= "000000000000";
      when "100011010011011" => color_data <= "010000110011";
      when "100011010011100" => color_data <= "011000100000";
      when "100011010011101" => color_data <= "011101000010";
      when "100011010011110" => color_data <= "011101000010";
      when "100011010011111" => color_data <= "011101000010";
      when "100011010100000" => color_data <= "011000100000";
      when "100011010100001" => color_data <= "101110010101";
      when "100011010100010" => color_data <= "111111111011";
      when "100011010100011" => color_data <= "111111101001";
      when "100011010100100" => color_data <= "111111101001";
      when "100011010100101" => color_data <= "111111101001";
      when "100011010100110" => color_data <= "111111101001";
      when "100011010100111" => color_data <= "111111101001";
      when "100011010101000" => color_data <= "111111101001";
      when "100011010101001" => color_data <= "111111101001";
      when "100011010101010" => color_data <= "111111101001";
      when "100011010101011" => color_data <= "111111101001";
      when "100011010101100" => color_data <= "111111101001";
      when "100011010101101" => color_data <= "111111101001";
      when "100011010101110" => color_data <= "111111101001";
      when "100011010101111" => color_data <= "111111101001";
      when "100011010110000" => color_data <= "111111101001";
      when "100011010110001" => color_data <= "111111101001";
      when "100011010110010" => color_data <= "111111101010";
      when "100011010110011" => color_data <= "111111111011";
      when "100011010110100" => color_data <= "111111101010";
      when "100011010110101" => color_data <= "111111101001";
      when "100011010110110" => color_data <= "111111101001";
      when "100011010110111" => color_data <= "111111101001";
      when "100011010111000" => color_data <= "111111101001";
      when "100011010111001" => color_data <= "111111101001";
      when "100011010111010" => color_data <= "111111101001";
      when "100011010111011" => color_data <= "111111101001";
      when "100011010111100" => color_data <= "111111101001";
      when "100011010111101" => color_data <= "111111101001";
      when "100011010111110" => color_data <= "111111101001";
      when "100011010111111" => color_data <= "111111101001";
      when "100011011000000" => color_data <= "111111101001";
      when "100011011000001" => color_data <= "111111101001";
      when "100011011000010" => color_data <= "111111111010";
      when "100011011000011" => color_data <= "110010110110";
      when "100011011000100" => color_data <= "011000100000";
      when "100011011000101" => color_data <= "011101000010";
      when "100011011000110" => color_data <= "011101000010";
      when "100011011000111" => color_data <= "011101000010";
      when "100011011001000" => color_data <= "011101000010";
      when "100011011001001" => color_data <= "011100110001";
      when "100011011001010" => color_data <= "011000110001";
      when "100011011001011" => color_data <= "000000000000";
      when "100011011001100" => color_data <= "000000000000";
      when "100011011001101" => color_data <= "000000000000";
      when "100011011001110" => color_data <= "000000000000";
      when "100011011001111" => color_data <= "000000000000";
      when "100011011010000" => color_data <= "000000000000";
      when "100011011010001" => color_data <= "000000000000";
      when "100011011010010" => color_data <= "000000000000";
      when "100011011010011" => color_data <= "000000000000";
      when "100011011010100" => color_data <= "000000000000";
      when "100011011010101" => color_data <= "000000000000";
      when "100011011010110" => color_data <= "000000000000";
      when "100011011010111" => color_data <= "000000000000";
      when "100011011011000" => color_data <= "000000000000";
      when "100011011011001" => color_data <= "000000000000";
      when "100011011011010" => color_data <= "000000000000";
      when "100011011011011" => color_data <= "000000000000";
      when "100011011011100" => color_data <= "000000000000";
      when "100011011011101" => color_data <= "000000000000";
      when "100011011011110" => color_data <= "000000000000";
      when "100011011011111" => color_data <= "000000000000";
      when "100011011100000" => color_data <= "000000000000";
      when "100011011100001" => color_data <= "000000000000";
      when "100011011100010" => color_data <= "000000000000";
      when "100011011100011" => color_data <= "000000000000";
      when "100011100000000" => color_data <= "000000000000";
      when "100011100000001" => color_data <= "000000000000";
      when "100011100000010" => color_data <= "000000000000";
      when "100011100000011" => color_data <= "000000000000";
      when "100011100000100" => color_data <= "000000000000";
      when "100011100000101" => color_data <= "000000000000";
      when "100011100000110" => color_data <= "000000000000";
      when "100011100000111" => color_data <= "000000000000";
      when "100011100001000" => color_data <= "000000000000";
      when "100011100001001" => color_data <= "000000000000";
      when "100011100001010" => color_data <= "000000000000";
      when "100011100001011" => color_data <= "000000000000";
      when "100011100001100" => color_data <= "000000000000";
      when "100011100001101" => color_data <= "000000000000";
      when "100011100001110" => color_data <= "000000000000";
      when "100011100001111" => color_data <= "000000000000";
      when "100011100010000" => color_data <= "000000000000";
      when "100011100010001" => color_data <= "000000000000";
      when "100011100010010" => color_data <= "000000000000";
      when "100011100010011" => color_data <= "000000000000";
      when "100011100010100" => color_data <= "000000000000";
      when "100011100010101" => color_data <= "000000000000";
      when "100011100010110" => color_data <= "000000000000";
      when "100011100010111" => color_data <= "000000000000";
      when "100011100011000" => color_data <= "000000000000";
      when "100011100011001" => color_data <= "000000000000";
      when "100011100011010" => color_data <= "000000000000";
      when "100011100011011" => color_data <= "010000110011";
      when "100011100011100" => color_data <= "011000100000";
      when "100011100011101" => color_data <= "011101000010";
      when "100011100011110" => color_data <= "011101000010";
      when "100011100011111" => color_data <= "011101000001";
      when "100011100100000" => color_data <= "010100100000";
      when "100011100100001" => color_data <= "101110010101";
      when "100011100100010" => color_data <= "111111111011";
      when "100011100100011" => color_data <= "111111101001";
      when "100011100100100" => color_data <= "111111101001";
      when "100011100100101" => color_data <= "111111101001";
      when "100011100100110" => color_data <= "111111101001";
      when "100011100100111" => color_data <= "111111101001";
      when "100011100101000" => color_data <= "111111101001";
      when "100011100101001" => color_data <= "111111101001";
      when "100011100101010" => color_data <= "111111101001";
      when "100011100101011" => color_data <= "111111101001";
      when "100011100101100" => color_data <= "111111101001";
      when "100011100101101" => color_data <= "111111101001";
      when "100011100101110" => color_data <= "111111101001";
      when "100011100101111" => color_data <= "111111101001";
      when "100011100110000" => color_data <= "111111101001";
      when "100011100110001" => color_data <= "111111101001";
      when "100011100110010" => color_data <= "111111101010";
      when "100011100110011" => color_data <= "111111111100";
      when "100011100110100" => color_data <= "111111101010";
      when "100011100110101" => color_data <= "111111101001";
      when "100011100110110" => color_data <= "111111101001";
      when "100011100110111" => color_data <= "111111101001";
      when "100011100111000" => color_data <= "111111101001";
      when "100011100111001" => color_data <= "111111101001";
      when "100011100111010" => color_data <= "111111101001";
      when "100011100111011" => color_data <= "111111101001";
      when "100011100111100" => color_data <= "111111101001";
      when "100011100111101" => color_data <= "111111101001";
      when "100011100111110" => color_data <= "111111101001";
      when "100011100111111" => color_data <= "111111101001";
      when "100011101000000" => color_data <= "111111101001";
      when "100011101000001" => color_data <= "111111101001";
      when "100011101000010" => color_data <= "111111111010";
      when "100011101000011" => color_data <= "110010110111";
      when "100011101000100" => color_data <= "011000100000";
      when "100011101000101" => color_data <= "011101000010";
      when "100011101000110" => color_data <= "011101000010";
      when "100011101000111" => color_data <= "011101000010";
      when "100011101001000" => color_data <= "011101000010";
      when "100011101001001" => color_data <= "011100110001";
      when "100011101001010" => color_data <= "011000110001";
      when "100011101001011" => color_data <= "000000000000";
      when "100011101001100" => color_data <= "000000000000";
      when "100011101001101" => color_data <= "000000000000";
      when "100011101001110" => color_data <= "000000000000";
      when "100011101001111" => color_data <= "000000000000";
      when "100011101010000" => color_data <= "000000000000";
      when "100011101010001" => color_data <= "000000000000";
      when "100011101010010" => color_data <= "000000000000";
      when "100011101010011" => color_data <= "000000000000";
      when "100011101010100" => color_data <= "000000000000";
      when "100011101010101" => color_data <= "000000000000";
      when "100011101010110" => color_data <= "000000000000";
      when "100011101010111" => color_data <= "000000000000";
      when "100011101011000" => color_data <= "000000000000";
      when "100011101011001" => color_data <= "000000000000";
      when "100011101011010" => color_data <= "000000000000";
      when "100011101011011" => color_data <= "000000000000";
      when "100011101011100" => color_data <= "000000000000";
      when "100011101011101" => color_data <= "000000000000";
      when "100011101011110" => color_data <= "000000000000";
      when "100011101011111" => color_data <= "000000000000";
      when "100011101100000" => color_data <= "000000000000";
      when "100011101100001" => color_data <= "000000000000";
      when "100011101100010" => color_data <= "000000000000";
      when "100011101100011" => color_data <= "000000000000";
      when "100011110000000" => color_data <= "000000000000";
      when "100011110000001" => color_data <= "000000000000";
      when "100011110000010" => color_data <= "000000000000";
      when "100011110000011" => color_data <= "000000000000";
      when "100011110000100" => color_data <= "000000000000";
      when "100011110000101" => color_data <= "000000000000";
      when "100011110000110" => color_data <= "000000000000";
      when "100011110000111" => color_data <= "000000000000";
      when "100011110001000" => color_data <= "000000000000";
      when "100011110001001" => color_data <= "000000000000";
      when "100011110001010" => color_data <= "000000000000";
      when "100011110001011" => color_data <= "000000000000";
      when "100011110001100" => color_data <= "000000000000";
      when "100011110001101" => color_data <= "000000000000";
      when "100011110001110" => color_data <= "000000000000";
      when "100011110001111" => color_data <= "000000000000";
      when "100011110010000" => color_data <= "000000000000";
      when "100011110010001" => color_data <= "000000000000";
      when "100011110010010" => color_data <= "000000000000";
      when "100011110010011" => color_data <= "000000000000";
      when "100011110010100" => color_data <= "000000000000";
      when "100011110010101" => color_data <= "000000000000";
      when "100011110010110" => color_data <= "000000000000";
      when "100011110010111" => color_data <= "000000000000";
      when "100011110011000" => color_data <= "000000000000";
      when "100011110011001" => color_data <= "000000000000";
      when "100011110011010" => color_data <= "000000000000";
      when "100011110011011" => color_data <= "010000110011";
      when "100011110011100" => color_data <= "011000100000";
      when "100011110011101" => color_data <= "011101000010";
      when "100011110011110" => color_data <= "011101000010";
      when "100011110011111" => color_data <= "011101000010";
      when "100011110100000" => color_data <= "010100100000";
      when "100011110100001" => color_data <= "101110010110";
      when "100011110100010" => color_data <= "111111111100";
      when "100011110100011" => color_data <= "111111111010";
      when "100011110100100" => color_data <= "111111111010";
      when "100011110100101" => color_data <= "111111111010";
      when "100011110100110" => color_data <= "111111111010";
      when "100011110100111" => color_data <= "111111111010";
      when "100011110101000" => color_data <= "111111111010";
      when "100011110101001" => color_data <= "111111111010";
      when "100011110101010" => color_data <= "111111111010";
      when "100011110101011" => color_data <= "111111111010";
      when "100011110101100" => color_data <= "111111111010";
      when "100011110101101" => color_data <= "111111111010";
      when "100011110101110" => color_data <= "111111111010";
      when "100011110101111" => color_data <= "111111111010";
      when "100011110110000" => color_data <= "111111111010";
      when "100011110110001" => color_data <= "111111111010";
      when "100011110110010" => color_data <= "111111111011";
      when "100011110110011" => color_data <= "111111111110";
      when "100011110110100" => color_data <= "111111111011";
      when "100011110110101" => color_data <= "111111111010";
      when "100011110110110" => color_data <= "111111111010";
      when "100011110110111" => color_data <= "111111111010";
      when "100011110111000" => color_data <= "111111111010";
      when "100011110111001" => color_data <= "111111111010";
      when "100011110111010" => color_data <= "111111111010";
      when "100011110111011" => color_data <= "111111111010";
      when "100011110111100" => color_data <= "111111111010";
      when "100011110111101" => color_data <= "111111111010";
      when "100011110111110" => color_data <= "111111111010";
      when "100011110111111" => color_data <= "111111111010";
      when "100011111000000" => color_data <= "111111111010";
      when "100011111000001" => color_data <= "111111111010";
      when "100011111000010" => color_data <= "111111111011";
      when "100011111000011" => color_data <= "110110110111";
      when "100011111000100" => color_data <= "011000100000";
      when "100011111000101" => color_data <= "011101000010";
      when "100011111000110" => color_data <= "011101000010";
      when "100011111000111" => color_data <= "011101000010";
      when "100011111001000" => color_data <= "011101000010";
      when "100011111001001" => color_data <= "011100110001";
      when "100011111001010" => color_data <= "011000110001";
      when "100011111001011" => color_data <= "000000000000";
      when "100011111001100" => color_data <= "000000000000";
      when "100011111001101" => color_data <= "000000000000";
      when "100011111001110" => color_data <= "000000000000";
      when "100011111001111" => color_data <= "000000000000";
      when "100011111010000" => color_data <= "000000000000";
      when "100011111010001" => color_data <= "000000000000";
      when "100011111010010" => color_data <= "000000000000";
      when "100011111010011" => color_data <= "000000000000";
      when "100011111010100" => color_data <= "000000000000";
      when "100011111010101" => color_data <= "000000000000";
      when "100011111010110" => color_data <= "000000000000";
      when "100011111010111" => color_data <= "000000000000";
      when "100011111011000" => color_data <= "000000000000";
      when "100011111011001" => color_data <= "000000000000";
      when "100011111011010" => color_data <= "000000000000";
      when "100011111011011" => color_data <= "000000000000";
      when "100011111011100" => color_data <= "000000000000";
      when "100011111011101" => color_data <= "000000000000";
      when "100011111011110" => color_data <= "000000000000";
      when "100011111011111" => color_data <= "000000000000";
      when "100011111100000" => color_data <= "000000000000";
      when "100011111100001" => color_data <= "000000000000";
      when "100011111100010" => color_data <= "000000000000";
      when "100011111100011" => color_data <= "000000000000";
      when "100100000000000" => color_data <= "000000000000";
      when "100100000000001" => color_data <= "000000000000";
      when "100100000000010" => color_data <= "000000000000";
      when "100100000000011" => color_data <= "000000000000";
      when "100100000000100" => color_data <= "000000000000";
      when "100100000000101" => color_data <= "000000000000";
      when "100100000000110" => color_data <= "000000000000";
      when "100100000000111" => color_data <= "000000000000";
      when "100100000001000" => color_data <= "000000000000";
      when "100100000001001" => color_data <= "000000000000";
      when "100100000001010" => color_data <= "000000000000";
      when "100100000001011" => color_data <= "000000000000";
      when "100100000001100" => color_data <= "000000000000";
      when "100100000001101" => color_data <= "000000000000";
      when "100100000001110" => color_data <= "000000000000";
      when "100100000001111" => color_data <= "000000000000";
      when "100100000010000" => color_data <= "000000000000";
      when "100100000010001" => color_data <= "000000000000";
      when "100100000010010" => color_data <= "000000000000";
      when "100100000010011" => color_data <= "000000000000";
      when "100100000010100" => color_data <= "000000000000";
      when "100100000010101" => color_data <= "000000000000";
      when "100100000010110" => color_data <= "000000000000";
      when "100100000010111" => color_data <= "000000000000";
      when "100100000011000" => color_data <= "000000000000";
      when "100100000011001" => color_data <= "000000000000";
      when "100100000011010" => color_data <= "000000000000";
      when "100100000011011" => color_data <= "010000110011";
      when "100100000011100" => color_data <= "010100000000";
      when "100100000011101" => color_data <= "011000110000";
      when "100100000011110" => color_data <= "011000110000";
      when "100100000011111" => color_data <= "011000110000";
      when "100100000100000" => color_data <= "011000100000";
      when "100100000100001" => color_data <= "011101000001";
      when "100100000100010" => color_data <= "100101110011";
      when "100100000100011" => color_data <= "100101100011";
      when "100100000100100" => color_data <= "100101100011";
      when "100100000100101" => color_data <= "100101100011";
      when "100100000100110" => color_data <= "100101100011";
      when "100100000100111" => color_data <= "100101100011";
      when "100100000101000" => color_data <= "100101100011";
      when "100100000101001" => color_data <= "100101100011";
      when "100100000101010" => color_data <= "100101100011";
      when "100100000101011" => color_data <= "100101100011";
      when "100100000101100" => color_data <= "100101100011";
      when "100100000101101" => color_data <= "100101100011";
      when "100100000101110" => color_data <= "100101100011";
      when "100100000101111" => color_data <= "100101100011";
      when "100100000110000" => color_data <= "100101100011";
      when "100100000110001" => color_data <= "100101100010";
      when "100100000110010" => color_data <= "100101100011";
      when "100100000110011" => color_data <= "100101110100";
      when "100100000110100" => color_data <= "100101100011";
      when "100100000110101" => color_data <= "100101100011";
      when "100100000110110" => color_data <= "100101100011";
      when "100100000110111" => color_data <= "100101100011";
      when "100100000111000" => color_data <= "100101100011";
      when "100100000111001" => color_data <= "100101100011";
      when "100100000111010" => color_data <= "100101100011";
      when "100100000111011" => color_data <= "100101100011";
      when "100100000111100" => color_data <= "100101100011";
      when "100100000111101" => color_data <= "100101100011";
      when "100100000111110" => color_data <= "100101100011";
      when "100100000111111" => color_data <= "100101100011";
      when "100100001000000" => color_data <= "100101100011";
      when "100100001000001" => color_data <= "100101100011";
      when "100100001000010" => color_data <= "100101110011";
      when "100100001000011" => color_data <= "100001010010";
      when "100100001000100" => color_data <= "011000100000";
      when "100100001000101" => color_data <= "011000110000";
      when "100100001000110" => color_data <= "011000110000";
      when "100100001000111" => color_data <= "011000110000";
      when "100100001001000" => color_data <= "011000110000";
      when "100100001001001" => color_data <= "011000100000";
      when "100100001001010" => color_data <= "010100100000";
      when "100100001001011" => color_data <= "000000000000";
      when "100100001001100" => color_data <= "000000000000";
      when "100100001001101" => color_data <= "000000000000";
      when "100100001001110" => color_data <= "000000000000";
      when "100100001001111" => color_data <= "000000000000";
      when "100100001010000" => color_data <= "000000000000";
      when "100100001010001" => color_data <= "000000000000";
      when "100100001010010" => color_data <= "000000000000";
      when "100100001010011" => color_data <= "000000000000";
      when "100100001010100" => color_data <= "000000000000";
      when "100100001010101" => color_data <= "000000000000";
      when "100100001010110" => color_data <= "000000000000";
      when "100100001010111" => color_data <= "000000000000";
      when "100100001011000" => color_data <= "000000000000";
      when "100100001011001" => color_data <= "000000000000";
      when "100100001011010" => color_data <= "000000000000";
      when "100100001011011" => color_data <= "000000000000";
      when "100100001011100" => color_data <= "000000000000";
      when "100100001011101" => color_data <= "000000000000";
      when "100100001011110" => color_data <= "000000000000";
      when "100100001011111" => color_data <= "000000000000";
      when "100100001100000" => color_data <= "000000000000";
      when "100100001100001" => color_data <= "000000000000";
      when "100100001100010" => color_data <= "000000000000";
      when "100100001100011" => color_data <= "000000000000";
      when "100100010000000" => color_data <= "000000000000";
      when "100100010000001" => color_data <= "000000000000";
      when "100100010000010" => color_data <= "000000000000";
      when "100100010000011" => color_data <= "000000000000";
      when "100100010000100" => color_data <= "000000000000";
      when "100100010000101" => color_data <= "000000000000";
      when "100100010000110" => color_data <= "000000000000";
      when "100100010000111" => color_data <= "000000000000";
      when "100100010001000" => color_data <= "000000000000";
      when "100100010001001" => color_data <= "000000000000";
      when "100100010001010" => color_data <= "000000000000";
      when "100100010001011" => color_data <= "000000000000";
      when "100100010001100" => color_data <= "000000000000";
      when "100100010001101" => color_data <= "000000000000";
      when "100100010001110" => color_data <= "000000000000";
      when "100100010001111" => color_data <= "000000000000";
      when "100100010010000" => color_data <= "000000000000";
      when "100100010010001" => color_data <= "000000000000";
      when "100100010010010" => color_data <= "000000000000";
      when "100100010010011" => color_data <= "000000000000";
      when "100100010010100" => color_data <= "000000000000";
      when "100100010010101" => color_data <= "000000000000";
      when "100100010010110" => color_data <= "000000000000";
      when "100100010010111" => color_data <= "000000000000";
      when "100100010011000" => color_data <= "000000000000";
      when "100100010011001" => color_data <= "000000000000";
      when "100100010011010" => color_data <= "000000000000";
      when "100100010011011" => color_data <= "001100110010";
      when "100100010011100" => color_data <= "010100110001";
      when "100100010011101" => color_data <= "010100110010";
      when "100100010011110" => color_data <= "010100110010";
      when "100100010011111" => color_data <= "010100110010";
      when "100100010100000" => color_data <= "010100110010";
      when "100100010100001" => color_data <= "010100110010";
      when "100100010100010" => color_data <= "010100100001";
      when "100100010100011" => color_data <= "010100110001";
      when "100100010100100" => color_data <= "010100110001";
      when "100100010100101" => color_data <= "010100110001";
      when "100100010100110" => color_data <= "010100110001";
      when "100100010100111" => color_data <= "010100110001";
      when "100100010101000" => color_data <= "010100110001";
      when "100100010101001" => color_data <= "010100110001";
      when "100100010101010" => color_data <= "010100110001";
      when "100100010101011" => color_data <= "010100110001";
      when "100100010101100" => color_data <= "010100110001";
      when "100100010101101" => color_data <= "010100110001";
      when "100100010101110" => color_data <= "010100110001";
      when "100100010101111" => color_data <= "010100110001";
      when "100100010110000" => color_data <= "010100110001";
      when "100100010110001" => color_data <= "010100110001";
      when "100100010110010" => color_data <= "010100110001";
      when "100100010110011" => color_data <= "010100100001";
      when "100100010110100" => color_data <= "010100110001";
      when "100100010110101" => color_data <= "010100110001";
      when "100100010110110" => color_data <= "010100110001";
      when "100100010110111" => color_data <= "010100110001";
      when "100100010111000" => color_data <= "010100110001";
      when "100100010111001" => color_data <= "010100110001";
      when "100100010111010" => color_data <= "010100110001";
      when "100100010111011" => color_data <= "010100110001";
      when "100100010111100" => color_data <= "010100110001";
      when "100100010111101" => color_data <= "010100110001";
      when "100100010111110" => color_data <= "010100110001";
      when "100100010111111" => color_data <= "010100110001";
      when "100100011000000" => color_data <= "010100110001";
      when "100100011000001" => color_data <= "010100110001";
      when "100100011000010" => color_data <= "010100100001";
      when "100100011000011" => color_data <= "010100110010";
      when "100100011000100" => color_data <= "010100110010";
      when "100100011000101" => color_data <= "010100110010";
      when "100100011000110" => color_data <= "010100110010";
      when "100100011000111" => color_data <= "010100110010";
      when "100100011001000" => color_data <= "010100110010";
      when "100100011001001" => color_data <= "010100110010";
      when "100100011001010" => color_data <= "010100110010";
      when "100100011001011" => color_data <= "000000000000";
      when "100100011001100" => color_data <= "000000000000";
      when "100100011001101" => color_data <= "000000000000";
      when "100100011001110" => color_data <= "000000000000";
      when "100100011001111" => color_data <= "000000000000";
      when "100100011010000" => color_data <= "000000000000";
      when "100100011010001" => color_data <= "000000000000";
      when "100100011010010" => color_data <= "000000000000";
      when "100100011010011" => color_data <= "000000000000";
      when "100100011010100" => color_data <= "000000000000";
      when "100100011010101" => color_data <= "000000000000";
      when "100100011010110" => color_data <= "000000000000";
      when "100100011010111" => color_data <= "000000000000";
      when "100100011011000" => color_data <= "000000000000";
      when "100100011011001" => color_data <= "000000000000";
      when "100100011011010" => color_data <= "000000000000";
      when "100100011011011" => color_data <= "000000000000";
      when "100100011011100" => color_data <= "000000000000";
      when "100100011011101" => color_data <= "000000000000";
      when "100100011011110" => color_data <= "000000000000";
      when "100100011011111" => color_data <= "000000000000";
      when "100100011100000" => color_data <= "000000000000";
      when "100100011100001" => color_data <= "000000000000";
      when "100100011100010" => color_data <= "000000000000";
      when "100100011100011" => color_data <= "000000000000";
      when "100100100000000" => color_data <= "000000000000";
      when "100100100000001" => color_data <= "000000000000";
      when "100100100000010" => color_data <= "000000000000";
      when "100100100000011" => color_data <= "000000000000";
      when "100100100000100" => color_data <= "000000000000";
      when "100100100000101" => color_data <= "000000000000";
      when "100100100000110" => color_data <= "000000000000";
      when "100100100000111" => color_data <= "000000000000";
      when "100100100001000" => color_data <= "000000000000";
      when "100100100001001" => color_data <= "000000000000";
      when "100100100001010" => color_data <= "000000000000";
      when "100100100001011" => color_data <= "000000000000";
      when "100100100001100" => color_data <= "000000000000";
      when "100100100001101" => color_data <= "000000000000";
      when "100100100001110" => color_data <= "000000000000";
      when "100100100001111" => color_data <= "000000000000";
      when "100100100010000" => color_data <= "000000000000";
      when "100100100010001" => color_data <= "000000000000";
      when "100100100010010" => color_data <= "000000000000";
      when "100100100010011" => color_data <= "000000000000";
      when "100100100010100" => color_data <= "000000000000";
      when "100100100010101" => color_data <= "000000000000";
      when "100100100010110" => color_data <= "000000000000";
      when "100100100010111" => color_data <= "000000000000";
      when "100100100011000" => color_data <= "000000000000";
      when "100100100011001" => color_data <= "000000000000";
      when "100100100011010" => color_data <= "000000000000";
      when "100100100011011" => color_data <= "000000000000";
      when "100100100011100" => color_data <= "000000000000";
      when "100100100011101" => color_data <= "000000000000";
      when "100100100011110" => color_data <= "000000000000";
      when "100100100011111" => color_data <= "000000000000";
      when "100100100100000" => color_data <= "000000000000";
      when "100100100100001" => color_data <= "000000000000";
      when "100100100100010" => color_data <= "000000000000";
      when "100100100100011" => color_data <= "000000000000";
      when "100100100100100" => color_data <= "000000000000";
      when "100100100100101" => color_data <= "000000000000";
      when "100100100100110" => color_data <= "000000000000";
      when "100100100100111" => color_data <= "000000000000";
      when "100100100101000" => color_data <= "000000000000";
      when "100100100101001" => color_data <= "000000000000";
      when "100100100101010" => color_data <= "000000000000";
      when "100100100101011" => color_data <= "000000000000";
      when "100100100101100" => color_data <= "000000000000";
      when "100100100101101" => color_data <= "000000000000";
      when "100100100101110" => color_data <= "000000000000";
      when "100100100101111" => color_data <= "000000000000";
      when "100100100110000" => color_data <= "000000000000";
      when "100100100110001" => color_data <= "000000000000";
      when "100100100110010" => color_data <= "000000000000";
      when "100100100110011" => color_data <= "000000000000";
      when "100100100110100" => color_data <= "000000000000";
      when "100100100110101" => color_data <= "000000000000";
      when "100100100110110" => color_data <= "000000000000";
      when "100100100110111" => color_data <= "000000000000";
      when "100100100111000" => color_data <= "000000000000";
      when "100100100111001" => color_data <= "000000000000";
      when "100100100111010" => color_data <= "000000000000";
      when "100100100111011" => color_data <= "000000000000";
      when "100100100111100" => color_data <= "000000000000";
      when "100100100111101" => color_data <= "000000000000";
      when "100100100111110" => color_data <= "000000000000";
      when "100100100111111" => color_data <= "000000000000";
      when "100100101000000" => color_data <= "000000000000";
      when "100100101000001" => color_data <= "000000000000";
      when "100100101000010" => color_data <= "000000000000";
      when "100100101000011" => color_data <= "000000000000";
      when "100100101000100" => color_data <= "000000000000";
      when "100100101000101" => color_data <= "000000000000";
      when "100100101000110" => color_data <= "000000000000";
      when "100100101000111" => color_data <= "000000000000";
      when "100100101001000" => color_data <= "000000000000";
      when "100100101001001" => color_data <= "000000000000";
      when "100100101001010" => color_data <= "000000000000";
      when "100100101001011" => color_data <= "000000000000";
      when "100100101001100" => color_data <= "000000000000";
      when "100100101001101" => color_data <= "000000000000";
      when "100100101001110" => color_data <= "000000000000";
      when "100100101001111" => color_data <= "000000000000";
      when "100100101010000" => color_data <= "000000000000";
      when "100100101010001" => color_data <= "000000000000";
      when "100100101010010" => color_data <= "000000000000";
      when "100100101010011" => color_data <= "000000000000";
      when "100100101010100" => color_data <= "000000000000";
      when "100100101010101" => color_data <= "000000000000";
      when "100100101010110" => color_data <= "000000000000";
      when "100100101010111" => color_data <= "000000000000";
      when "100100101011000" => color_data <= "000000000000";
      when "100100101011001" => color_data <= "000000000000";
      when "100100101011010" => color_data <= "000000000000";
      when "100100101011011" => color_data <= "000000000000";
      when "100100101011100" => color_data <= "000000000000";
      when "100100101011101" => color_data <= "000000000000";
      when "100100101011110" => color_data <= "000000000000";
      when "100100101011111" => color_data <= "000000000000";
      when "100100101100000" => color_data <= "000000000000";
      when "100100101100001" => color_data <= "000000000000";
      when "100100101100010" => color_data <= "000000000000";
      when "100100101100011" => color_data <= "000000000000";
      when "100100110000000" => color_data <= "000000000000";
      when "100100110000001" => color_data <= "000000000000";
      when "100100110000010" => color_data <= "000000000000";
      when "100100110000011" => color_data <= "000000000000";
      when "100100110000100" => color_data <= "000000000000";
      when "100100110000101" => color_data <= "000000000000";
      when "100100110000110" => color_data <= "000000000000";
      when "100100110000111" => color_data <= "000000000000";
      when "100100110001000" => color_data <= "000000000000";
      when "100100110001001" => color_data <= "000000000000";
      when "100100110001010" => color_data <= "000000000000";
      when "100100110001011" => color_data <= "000000000000";
      when "100100110001100" => color_data <= "000000000000";
      when "100100110001101" => color_data <= "000000000000";
      when "100100110001110" => color_data <= "000000000000";
      when "100100110001111" => color_data <= "000000000000";
      when "100100110010000" => color_data <= "000000000000";
      when "100100110010001" => color_data <= "000000000000";
      when "100100110010010" => color_data <= "000000000000";
      when "100100110010011" => color_data <= "000000000000";
      when "100100110010100" => color_data <= "000000000000";
      when "100100110010101" => color_data <= "000000000000";
      when "100100110010110" => color_data <= "000000000000";
      when "100100110010111" => color_data <= "000000000000";
      when "100100110011000" => color_data <= "000000000000";
      when "100100110011001" => color_data <= "000000000000";
      when "100100110011010" => color_data <= "000000000000";
      when "100100110011011" => color_data <= "000000000000";
      when "100100110011100" => color_data <= "000000000000";
      when "100100110011101" => color_data <= "000000000000";
      when "100100110011110" => color_data <= "000000000000";
      when "100100110011111" => color_data <= "000000000000";
      when "100100110100000" => color_data <= "000000000000";
      when "100100110100001" => color_data <= "000000000000";
      when "100100110100010" => color_data <= "000000000000";
      when "100100110100011" => color_data <= "000000000000";
      when "100100110100100" => color_data <= "000000000000";
      when "100100110100101" => color_data <= "000000000000";
      when "100100110100110" => color_data <= "000000000000";
      when "100100110100111" => color_data <= "000000000000";
      when "100100110101000" => color_data <= "000000000000";
      when "100100110101001" => color_data <= "000000000000";
      when "100100110101010" => color_data <= "000000000000";
      when "100100110101011" => color_data <= "000000000000";
      when "100100110101100" => color_data <= "000000000000";
      when "100100110101101" => color_data <= "000000000000";
      when "100100110101110" => color_data <= "000000000000";
      when "100100110101111" => color_data <= "000000000000";
      when "100100110110000" => color_data <= "000000000000";
      when "100100110110001" => color_data <= "000000000000";
      when "100100110110010" => color_data <= "000000000000";
      when "100100110110011" => color_data <= "000000000000";
      when "100100110110100" => color_data <= "000000000000";
      when "100100110110101" => color_data <= "000000000000";
      when "100100110110110" => color_data <= "000000000000";
      when "100100110110111" => color_data <= "000000000000";
      when "100100110111000" => color_data <= "000000000000";
      when "100100110111001" => color_data <= "000000000000";
      when "100100110111010" => color_data <= "000000000000";
      when "100100110111011" => color_data <= "000000000000";
      when "100100110111100" => color_data <= "000000000000";
      when "100100110111101" => color_data <= "000000000000";
      when "100100110111110" => color_data <= "000000000000";
      when "100100110111111" => color_data <= "000000000000";
      when "100100111000000" => color_data <= "000000000000";
      when "100100111000001" => color_data <= "000000000000";
      when "100100111000010" => color_data <= "000000000000";
      when "100100111000011" => color_data <= "000000000000";
      when "100100111000100" => color_data <= "000000000000";
      when "100100111000101" => color_data <= "000000000000";
      when "100100111000110" => color_data <= "000000000000";
      when "100100111000111" => color_data <= "000000000000";
      when "100100111001000" => color_data <= "000000000000";
      when "100100111001001" => color_data <= "000000000000";
      when "100100111001010" => color_data <= "000000000000";
      when "100100111001011" => color_data <= "000000000000";
      when "100100111001100" => color_data <= "000000000000";
      when "100100111001101" => color_data <= "000000000000";
      when "100100111001110" => color_data <= "000000000000";
      when "100100111001111" => color_data <= "000000000000";
      when "100100111010000" => color_data <= "000000000000";
      when "100100111010001" => color_data <= "000000000000";
      when "100100111010010" => color_data <= "000000000000";
      when "100100111010011" => color_data <= "000000000000";
      when "100100111010100" => color_data <= "000000000000";
      when "100100111010101" => color_data <= "000000000000";
      when "100100111010110" => color_data <= "000000000000";
      when "100100111010111" => color_data <= "000000000000";
      when "100100111011000" => color_data <= "000000000000";
      when "100100111011001" => color_data <= "000000000000";
      when "100100111011010" => color_data <= "000000000000";
      when "100100111011011" => color_data <= "000000000000";
      when "100100111011100" => color_data <= "000000000000";
      when "100100111011101" => color_data <= "000000000000";
      when "100100111011110" => color_data <= "000000000000";
      when "100100111011111" => color_data <= "000000000000";
      when "100100111100000" => color_data <= "000000000000";
      when "100100111100001" => color_data <= "000000000000";
      when "100100111100010" => color_data <= "000000000000";
      when "100100111100011" => color_data <= "000000000000";
      when "100101000000000" => color_data <= "000000000000";
      when "100101000000001" => color_data <= "000000000000";
      when "100101000000010" => color_data <= "000000000000";
      when "100101000000011" => color_data <= "000000000000";
      when "100101000000100" => color_data <= "000000000000";
      when "100101000000101" => color_data <= "000000000000";
      when "100101000000110" => color_data <= "000000000000";
      when "100101000000111" => color_data <= "000000000000";
      when "100101000001000" => color_data <= "000000000000";
      when "100101000001001" => color_data <= "000000000000";
      when "100101000001010" => color_data <= "000000000000";
      when "100101000001011" => color_data <= "000000000000";
      when "100101000001100" => color_data <= "000000000000";
      when "100101000001101" => color_data <= "000000000000";
      when "100101000001110" => color_data <= "000000000000";
      when "100101000001111" => color_data <= "000000000000";
      when "100101000010000" => color_data <= "000000000000";
      when "100101000010001" => color_data <= "000000000000";
      when "100101000010010" => color_data <= "000000000000";
      when "100101000010011" => color_data <= "000000000000";
      when "100101000010100" => color_data <= "000000000000";
      when "100101000010101" => color_data <= "000000000000";
      when "100101000010110" => color_data <= "000000000000";
      when "100101000010111" => color_data <= "000000000000";
      when "100101000011000" => color_data <= "000000000000";
      when "100101000011001" => color_data <= "000000000000";
      when "100101000011010" => color_data <= "000000000000";
      when "100101000011011" => color_data <= "000000000000";
      when "100101000011100" => color_data <= "000000000000";
      when "100101000011101" => color_data <= "000000000000";
      when "100101000011110" => color_data <= "000000000000";
      when "100101000011111" => color_data <= "000000000000";
      when "100101000100000" => color_data <= "000000000000";
      when "100101000100001" => color_data <= "000000000000";
      when "100101000100010" => color_data <= "000000000000";
      when "100101000100011" => color_data <= "000000000000";
      when "100101000100100" => color_data <= "000000000000";
      when "100101000100101" => color_data <= "000000000000";
      when "100101000100110" => color_data <= "000000000000";
      when "100101000100111" => color_data <= "000000000000";
      when "100101000101000" => color_data <= "000000000000";
      when "100101000101001" => color_data <= "000000000000";
      when "100101000101010" => color_data <= "000000000000";
      when "100101000101011" => color_data <= "000000000000";
      when "100101000101100" => color_data <= "000000000000";
      when "100101000101101" => color_data <= "000000000000";
      when "100101000101110" => color_data <= "000000000000";
      when "100101000101111" => color_data <= "000000000000";
      when "100101000110000" => color_data <= "000000000000";
      when "100101000110001" => color_data <= "000000000000";
      when "100101000110010" => color_data <= "000000000000";
      when "100101000110011" => color_data <= "000000000000";
      when "100101000110100" => color_data <= "000000000000";
      when "100101000110101" => color_data <= "000000000000";
      when "100101000110110" => color_data <= "000000000000";
      when "100101000110111" => color_data <= "000000000000";
      when "100101000111000" => color_data <= "000000000000";
      when "100101000111001" => color_data <= "000000000000";
      when "100101000111010" => color_data <= "000000000000";
      when "100101000111011" => color_data <= "000000000000";
      when "100101000111100" => color_data <= "000000000000";
      when "100101000111101" => color_data <= "000000000000";
      when "100101000111110" => color_data <= "000000000000";
      when "100101000111111" => color_data <= "000000000000";
      when "100101001000000" => color_data <= "000000000000";
      when "100101001000001" => color_data <= "000000000000";
      when "100101001000010" => color_data <= "000000000000";
      when "100101001000011" => color_data <= "000000000000";
      when "100101001000100" => color_data <= "000000000000";
      when "100101001000101" => color_data <= "000000000000";
      when "100101001000110" => color_data <= "000000000000";
      when "100101001000111" => color_data <= "000000000000";
      when "100101001001000" => color_data <= "000000000000";
      when "100101001001001" => color_data <= "000000000000";
      when "100101001001010" => color_data <= "000000000000";
      when "100101001001011" => color_data <= "000000000000";
      when "100101001001100" => color_data <= "000000000000";
      when "100101001001101" => color_data <= "000000000000";
      when "100101001001110" => color_data <= "000000000000";
      when "100101001001111" => color_data <= "000000000000";
      when "100101001010000" => color_data <= "000000000000";
      when "100101001010001" => color_data <= "000000000000";
      when "100101001010010" => color_data <= "000000000000";
      when "100101001010011" => color_data <= "000000000000";
      when "100101001010100" => color_data <= "000000000000";
      when "100101001010101" => color_data <= "000000000000";
      when "100101001010110" => color_data <= "000000000000";
      when "100101001010111" => color_data <= "000000000000";
      when "100101001011000" => color_data <= "000000000000";
      when "100101001011001" => color_data <= "000000000000";
      when "100101001011010" => color_data <= "000000000000";
      when "100101001011011" => color_data <= "000000000000";
      when "100101001011100" => color_data <= "000000000000";
      when "100101001011101" => color_data <= "000000000000";
      when "100101001011110" => color_data <= "000000000000";
      when "100101001011111" => color_data <= "000000000000";
      when "100101001100000" => color_data <= "000000000000";
      when "100101001100001" => color_data <= "000000000000";
      when "100101001100010" => color_data <= "000000000000";
      when "100101001100011" => color_data <= "000000000000";
      when others => color_data <= (others => '0');
    end case;
  end process;
end Behavioral;
