library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity brick_rom is
  Port (
    clk        : in  std_logic;
    row        : in  std_logic_vector(9 downto 0);
    col        : in  std_logic_vector(9 downto 0);
    color_data : out std_logic_vector(11 downto 0)
  );
end entity;

architecture Behavioral of brick_rom is
  signal addr : std_logic_vector(10 downto 0);
  signal row_reg : std_logic_vector(4 downto 0);
  signal col_reg : std_logic_vector(5 downto 0);
begin

  process(clk)
  begin
    if rising_edge(clk) then
      row_reg <= row(4 downto 0);
      col_reg <= col(5 downto 0);
    end if;
  end process;

  addr <= row_reg & col_reg;

  process(addr)
  begin
    case addr is
      when "00000000000" => color_data <= "110001100011";
      when "00000000001" => color_data <= "110001000010";
      when "00000000010" => color_data <= "110001010010";
      when "00000000011" => color_data <= "110001010010";
      when "00000000100" => color_data <= "011101000010";
      when "00000000101" => color_data <= "100101000010";
      when "00000000110" => color_data <= "110101010010";
      when "00000000111" => color_data <= "110001010010";
      when "00000001000" => color_data <= "110001010010";
      when "00000001001" => color_data <= "110001010010";
      when "00000001010" => color_data <= "110001010010";
      when "00000001011" => color_data <= "110001010010";
      when "00000001100" => color_data <= "110001010010";
      when "00000001101" => color_data <= "110001010010";
      when "00000001110" => color_data <= "110001010010";
      when "00000001111" => color_data <= "110001010010";
      when "00000010000" => color_data <= "110001010010";
      when "00000010001" => color_data <= "110001010010";
      when "00000010010" => color_data <= "110001010010";
      when "00000010011" => color_data <= "110001010010";
      when "00000010100" => color_data <= "110001010010";
      when "00000010101" => color_data <= "110001010010";
      when "00000010110" => color_data <= "101101010010";
      when "00000010111" => color_data <= "011101000010";
      when "00000011000" => color_data <= "101101010010";
      when "00000011001" => color_data <= "110001010010";
      when "00000011010" => color_data <= "110001010010";
      when "00000011011" => color_data <= "110001010010";
      when "00000011100" => color_data <= "110001010010";
      when "00000011101" => color_data <= "110001010010";
      when "00000011110" => color_data <= "110001010010";
      when "00000011111" => color_data <= "110001010010";
      when "00000100000" => color_data <= "110001010010";
      when "00000100001" => color_data <= "110001010010";
      when "00000100010" => color_data <= "110001010010";
      when "00000100011" => color_data <= "110001010010";
      when "00000100100" => color_data <= "110001010010";
      when "00000100101" => color_data <= "110001010010";
      when "00000100110" => color_data <= "110001010010";
      when "00000100111" => color_data <= "110001010010";
      when "00000101000" => color_data <= "110101010010";
      when "00000101001" => color_data <= "100001000010";
      when "00000101010" => color_data <= "011101000010";
      when "00000101011" => color_data <= "110001010010";
      when "00000101100" => color_data <= "110001010010";
      when "00000101101" => color_data <= "110001010010";
      when "00000101110" => color_data <= "110001010010";
      when "00000101111" => color_data <= "110001010010";
      when "00000110000" => color_data <= "110001010010";
      when "00000110001" => color_data <= "110001010010";
      when "00000110010" => color_data <= "110001010010";
      when "00000110011" => color_data <= "110001010010";
      when "00000110100" => color_data <= "110001010010";
      when "00000110101" => color_data <= "110001010010";
      when "00000110110" => color_data <= "110001010010";
      when "00000110111" => color_data <= "110001010010";
      when "00000111000" => color_data <= "110001010010";
      when "00000111001" => color_data <= "110001010010";
      when "00000111010" => color_data <= "110001010010";
      when "00000111011" => color_data <= "110101010010";
      when "00000111100" => color_data <= "100001000010";
      when "00000111101" => color_data <= "100101000010";
      when "00000111110" => color_data <= "110101010010";
      when "00000111111" => color_data <= "110001100011";
      when "00001000000" => color_data <= "110001010010";
      when "00001000001" => color_data <= "110001000010";
      when "00001000010" => color_data <= "110001000010";
      when "00001000011" => color_data <= "110001010010";
      when "00001000100" => color_data <= "011000110010";
      when "00001000101" => color_data <= "100101000010";
      when "00001000110" => color_data <= "110101010010";
      when "00001000111" => color_data <= "110001000010";
      when "00001001000" => color_data <= "110001000010";
      when "00001001001" => color_data <= "110001000010";
      when "00001001010" => color_data <= "110001000010";
      when "00001001011" => color_data <= "110001000010";
      when "00001001100" => color_data <= "110001000010";
      when "00001001101" => color_data <= "110001000010";
      when "00001001110" => color_data <= "110001000010";
      when "00001001111" => color_data <= "110001000010";
      when "00001010000" => color_data <= "110001000010";
      when "00001010001" => color_data <= "110001000010";
      when "00001010010" => color_data <= "110001000010";
      when "00001010011" => color_data <= "110001000010";
      when "00001010100" => color_data <= "110001000010";
      when "00001010101" => color_data <= "110001010010";
      when "00001010110" => color_data <= "101101000010";
      when "00001010111" => color_data <= "011000110010";
      when "00001011000" => color_data <= "101101000010";
      when "00001011001" => color_data <= "110001010010";
      when "00001011010" => color_data <= "110001000010";
      when "00001011011" => color_data <= "110001000010";
      when "00001011100" => color_data <= "110001000010";
      when "00001011101" => color_data <= "110001000010";
      when "00001011110" => color_data <= "110001000010";
      when "00001011111" => color_data <= "110001000010";
      when "00001100000" => color_data <= "110001000010";
      when "00001100001" => color_data <= "110001000010";
      when "00001100010" => color_data <= "110001000010";
      when "00001100011" => color_data <= "110001000010";
      when "00001100100" => color_data <= "110001000010";
      when "00001100101" => color_data <= "110001000010";
      when "00001100110" => color_data <= "110001000010";
      when "00001100111" => color_data <= "110001000010";
      when "00001101000" => color_data <= "110101010010";
      when "00001101001" => color_data <= "100001000010";
      when "00001101010" => color_data <= "011000110010";
      when "00001101011" => color_data <= "110001010010";
      when "00001101100" => color_data <= "110001010010";
      when "00001101101" => color_data <= "110001000010";
      when "00001101110" => color_data <= "110001000010";
      when "00001101111" => color_data <= "110001000010";
      when "00001110000" => color_data <= "110001000010";
      when "00001110001" => color_data <= "110001000010";
      when "00001110010" => color_data <= "110001000010";
      when "00001110011" => color_data <= "110001000010";
      when "00001110100" => color_data <= "110001000010";
      when "00001110101" => color_data <= "110001000010";
      when "00001110110" => color_data <= "110001000010";
      when "00001110111" => color_data <= "110001000010";
      when "00001111000" => color_data <= "110001000010";
      when "00001111001" => color_data <= "110001000010";
      when "00001111010" => color_data <= "110001000010";
      when "00001111011" => color_data <= "110001010010";
      when "00001111100" => color_data <= "011100110010";
      when "00001111101" => color_data <= "100101000010";
      when "00001111110" => color_data <= "110101010010";
      when "00001111111" => color_data <= "110001010010";
      when "00010000000" => color_data <= "110001010010";
      when "00010000001" => color_data <= "110001000010";
      when "00010000010" => color_data <= "110001000010";
      when "00010000011" => color_data <= "110001010010";
      when "00010000100" => color_data <= "011000110010";
      when "00010000101" => color_data <= "100101000010";
      when "00010000110" => color_data <= "110101010010";
      when "00010000111" => color_data <= "110001000010";
      when "00010001000" => color_data <= "110001000010";
      when "00010001001" => color_data <= "110001000010";
      when "00010001010" => color_data <= "110001000010";
      when "00010001011" => color_data <= "110001000010";
      when "00010001100" => color_data <= "110001000010";
      when "00010001101" => color_data <= "110001000010";
      when "00010001110" => color_data <= "110001000010";
      when "00010001111" => color_data <= "110001000010";
      when "00010010000" => color_data <= "110001000010";
      when "00010010001" => color_data <= "110001000010";
      when "00010010010" => color_data <= "110001000010";
      when "00010010011" => color_data <= "110001000010";
      when "00010010100" => color_data <= "110001000010";
      when "00010010101" => color_data <= "110001010010";
      when "00010010110" => color_data <= "101101000010";
      when "00010010111" => color_data <= "011000110010";
      when "00010011000" => color_data <= "101101000010";
      when "00010011001" => color_data <= "110001010010";
      when "00010011010" => color_data <= "110001000010";
      when "00010011011" => color_data <= "110001000010";
      when "00010011100" => color_data <= "110001000010";
      when "00010011101" => color_data <= "110001000010";
      when "00010011110" => color_data <= "110001000010";
      when "00010011111" => color_data <= "110001000010";
      when "00010100000" => color_data <= "110001000010";
      when "00010100001" => color_data <= "110001000010";
      when "00010100010" => color_data <= "110001000010";
      when "00010100011" => color_data <= "110001000010";
      when "00010100100" => color_data <= "110001000010";
      when "00010100101" => color_data <= "110001000010";
      when "00010100110" => color_data <= "110001000010";
      when "00010100111" => color_data <= "110001000010";
      when "00010101000" => color_data <= "110101010010";
      when "00010101001" => color_data <= "100001000010";
      when "00010101010" => color_data <= "011000110010";
      when "00010101011" => color_data <= "110001010010";
      when "00010101100" => color_data <= "110001010010";
      when "00010101101" => color_data <= "110001000010";
      when "00010101110" => color_data <= "110001000010";
      when "00010101111" => color_data <= "110001000010";
      when "00010110000" => color_data <= "110001000010";
      when "00010110001" => color_data <= "110001000010";
      when "00010110010" => color_data <= "110001000010";
      when "00010110011" => color_data <= "110001000010";
      when "00010110100" => color_data <= "110001000010";
      when "00010110101" => color_data <= "110001000010";
      when "00010110110" => color_data <= "110001000010";
      when "00010110111" => color_data <= "110001000010";
      when "00010111000" => color_data <= "110001000010";
      when "00010111001" => color_data <= "110001000010";
      when "00010111010" => color_data <= "110001000010";
      when "00010111011" => color_data <= "110001010010";
      when "00010111100" => color_data <= "011100110010";
      when "00010111101" => color_data <= "100101000010";
      when "00010111110" => color_data <= "110101010010";
      when "00010111111" => color_data <= "110001010010";
      when "00011000000" => color_data <= "110001010010";
      when "00011000001" => color_data <= "110001000010";
      when "00011000010" => color_data <= "110001000010";
      when "00011000011" => color_data <= "110001010010";
      when "00011000100" => color_data <= "011000110010";
      when "00011000101" => color_data <= "100101000010";
      when "00011000110" => color_data <= "110101010010";
      when "00011000111" => color_data <= "110001000010";
      when "00011001000" => color_data <= "110001000010";
      when "00011001001" => color_data <= "110001000010";
      when "00011001010" => color_data <= "110001000010";
      when "00011001011" => color_data <= "110001000010";
      when "00011001100" => color_data <= "110001000010";
      when "00011001101" => color_data <= "110001000010";
      when "00011001110" => color_data <= "110001000010";
      when "00011001111" => color_data <= "110001000010";
      when "00011010000" => color_data <= "110001000010";
      when "00011010001" => color_data <= "110001000010";
      when "00011010010" => color_data <= "110001000010";
      when "00011010011" => color_data <= "110001000010";
      when "00011010100" => color_data <= "110001000010";
      when "00011010101" => color_data <= "110001010010";
      when "00011010110" => color_data <= "101101000010";
      when "00011010111" => color_data <= "011000110010";
      when "00011011000" => color_data <= "101101000010";
      when "00011011001" => color_data <= "110001010010";
      when "00011011010" => color_data <= "110001000010";
      when "00011011011" => color_data <= "110001000010";
      when "00011011100" => color_data <= "110001000010";
      when "00011011101" => color_data <= "110001000010";
      when "00011011110" => color_data <= "110001000010";
      when "00011011111" => color_data <= "110001000010";
      when "00011100000" => color_data <= "110001000010";
      when "00011100001" => color_data <= "110001000010";
      when "00011100010" => color_data <= "110001000010";
      when "00011100011" => color_data <= "110001000010";
      when "00011100100" => color_data <= "110001000010";
      when "00011100101" => color_data <= "110001000010";
      when "00011100110" => color_data <= "110001000010";
      when "00011100111" => color_data <= "110001000010";
      when "00011101000" => color_data <= "110101010010";
      when "00011101001" => color_data <= "100001000010";
      when "00011101010" => color_data <= "011000110010";
      when "00011101011" => color_data <= "110001010010";
      when "00011101100" => color_data <= "110001010010";
      when "00011101101" => color_data <= "110001000010";
      when "00011101110" => color_data <= "110001000010";
      when "00011101111" => color_data <= "110001000010";
      when "00011110000" => color_data <= "110001000010";
      when "00011110001" => color_data <= "110001000010";
      when "00011110010" => color_data <= "110001000010";
      when "00011110011" => color_data <= "110001000010";
      when "00011110100" => color_data <= "110001000010";
      when "00011110101" => color_data <= "110001000010";
      when "00011110110" => color_data <= "110001000010";
      when "00011110111" => color_data <= "110001000010";
      when "00011111000" => color_data <= "110001000010";
      when "00011111001" => color_data <= "110001000010";
      when "00011111010" => color_data <= "110001000010";
      when "00011111011" => color_data <= "110001010010";
      when "00011111100" => color_data <= "011100110010";
      when "00011111101" => color_data <= "100101000010";
      when "00011111110" => color_data <= "110101010010";
      when "00011111111" => color_data <= "110001010010";
      when "00100000000" => color_data <= "110001010010";
      when "00100000001" => color_data <= "110001000010";
      when "00100000010" => color_data <= "110001000010";
      when "00100000011" => color_data <= "110001010010";
      when "00100000100" => color_data <= "011000110010";
      when "00100000101" => color_data <= "100101000010";
      when "00100000110" => color_data <= "110101010010";
      when "00100000111" => color_data <= "110001000010";
      when "00100001000" => color_data <= "110001000010";
      when "00100001001" => color_data <= "110001000010";
      when "00100001010" => color_data <= "110001000010";
      when "00100001011" => color_data <= "110001000010";
      when "00100001100" => color_data <= "110001000010";
      when "00100001101" => color_data <= "110001000010";
      when "00100001110" => color_data <= "110001000010";
      when "00100001111" => color_data <= "110001000010";
      when "00100010000" => color_data <= "110001000010";
      when "00100010001" => color_data <= "110001000010";
      when "00100010010" => color_data <= "110001000010";
      when "00100010011" => color_data <= "110001000010";
      when "00100010100" => color_data <= "110001000010";
      when "00100010101" => color_data <= "110001010010";
      when "00100010110" => color_data <= "101101000010";
      when "00100010111" => color_data <= "011000110010";
      when "00100011000" => color_data <= "101101000010";
      when "00100011001" => color_data <= "110001010010";
      when "00100011010" => color_data <= "110001000010";
      when "00100011011" => color_data <= "110001000010";
      when "00100011100" => color_data <= "110001000010";
      when "00100011101" => color_data <= "110001000010";
      when "00100011110" => color_data <= "110001000010";
      when "00100011111" => color_data <= "110001000010";
      when "00100100000" => color_data <= "110001000010";
      when "00100100001" => color_data <= "110001000010";
      when "00100100010" => color_data <= "110001000010";
      when "00100100011" => color_data <= "110001000010";
      when "00100100100" => color_data <= "110001000010";
      when "00100100101" => color_data <= "110001000010";
      when "00100100110" => color_data <= "110001000010";
      when "00100100111" => color_data <= "110001000010";
      when "00100101000" => color_data <= "110101010010";
      when "00100101001" => color_data <= "100001000010";
      when "00100101010" => color_data <= "011000110010";
      when "00100101011" => color_data <= "110001010010";
      when "00100101100" => color_data <= "110001010010";
      when "00100101101" => color_data <= "110001000010";
      when "00100101110" => color_data <= "110001000010";
      when "00100101111" => color_data <= "110001000010";
      when "00100110000" => color_data <= "110001000010";
      when "00100110001" => color_data <= "110001000010";
      when "00100110010" => color_data <= "110001000010";
      when "00100110011" => color_data <= "110001000010";
      when "00100110100" => color_data <= "110001000010";
      when "00100110101" => color_data <= "110001000010";
      when "00100110110" => color_data <= "110001000010";
      when "00100110111" => color_data <= "110001000010";
      when "00100111000" => color_data <= "110001000010";
      when "00100111001" => color_data <= "110001000010";
      when "00100111010" => color_data <= "110001000010";
      when "00100111011" => color_data <= "110001010010";
      when "00100111100" => color_data <= "011100110010";
      when "00100111101" => color_data <= "100101000010";
      when "00100111110" => color_data <= "110101010010";
      when "00100111111" => color_data <= "110001010010";
      when "00101000000" => color_data <= "110001010010";
      when "00101000001" => color_data <= "110001000010";
      when "00101000010" => color_data <= "110001000010";
      when "00101000011" => color_data <= "110001010010";
      when "00101000100" => color_data <= "011000110010";
      when "00101000101" => color_data <= "100101000010";
      when "00101000110" => color_data <= "110101010010";
      when "00101000111" => color_data <= "110001000010";
      when "00101001000" => color_data <= "110001000010";
      when "00101001001" => color_data <= "110001000010";
      when "00101001010" => color_data <= "110001000010";
      when "00101001011" => color_data <= "110001000010";
      when "00101001100" => color_data <= "110001000010";
      when "00101001101" => color_data <= "110001000010";
      when "00101001110" => color_data <= "110001000010";
      when "00101001111" => color_data <= "110001000010";
      when "00101010000" => color_data <= "110001000010";
      when "00101010001" => color_data <= "110001000010";
      when "00101010010" => color_data <= "110001000010";
      when "00101010011" => color_data <= "110001000010";
      when "00101010100" => color_data <= "110001000010";
      when "00101010101" => color_data <= "110001010010";
      when "00101010110" => color_data <= "101101000010";
      when "00101010111" => color_data <= "011000110010";
      when "00101011000" => color_data <= "101101000010";
      when "00101011001" => color_data <= "110001010010";
      when "00101011010" => color_data <= "110001000010";
      when "00101011011" => color_data <= "110001000010";
      when "00101011100" => color_data <= "110001000010";
      when "00101011101" => color_data <= "110001000010";
      when "00101011110" => color_data <= "110001000010";
      when "00101011111" => color_data <= "110001000010";
      when "00101100000" => color_data <= "110001000010";
      when "00101100001" => color_data <= "110001000010";
      when "00101100010" => color_data <= "110001000010";
      when "00101100011" => color_data <= "110001000010";
      when "00101100100" => color_data <= "110001000010";
      when "00101100101" => color_data <= "110001000010";
      when "00101100110" => color_data <= "110001000010";
      when "00101100111" => color_data <= "110001000010";
      when "00101101000" => color_data <= "110101010010";
      when "00101101001" => color_data <= "100001000010";
      when "00101101010" => color_data <= "011000110010";
      when "00101101011" => color_data <= "110001010010";
      when "00101101100" => color_data <= "110001010010";
      when "00101101101" => color_data <= "110001000010";
      when "00101101110" => color_data <= "110001000010";
      when "00101101111" => color_data <= "110001000010";
      when "00101110000" => color_data <= "110001000010";
      when "00101110001" => color_data <= "110001000010";
      when "00101110010" => color_data <= "110001000010";
      when "00101110011" => color_data <= "110001000010";
      when "00101110100" => color_data <= "110001000010";
      when "00101110101" => color_data <= "110001000010";
      when "00101110110" => color_data <= "110001000010";
      when "00101110111" => color_data <= "110001000010";
      when "00101111000" => color_data <= "110001000010";
      when "00101111001" => color_data <= "110001000010";
      when "00101111010" => color_data <= "110001000010";
      when "00101111011" => color_data <= "110101010010";
      when "00101111100" => color_data <= "011100110010";
      when "00101111101" => color_data <= "100101000010";
      when "00101111110" => color_data <= "110101010010";
      when "00101111111" => color_data <= "110001010010";
      when "00110000000" => color_data <= "110001010010";
      when "00110000001" => color_data <= "110001010010";
      when "00110000010" => color_data <= "110001010010";
      when "00110000011" => color_data <= "110101010010";
      when "00110000100" => color_data <= "011000110010";
      when "00110000101" => color_data <= "100101000010";
      when "00110000110" => color_data <= "110101010010";
      when "00110000111" => color_data <= "110001010010";
      when "00110001000" => color_data <= "110001010010";
      when "00110001001" => color_data <= "110001010010";
      when "00110001010" => color_data <= "110001010010";
      when "00110001011" => color_data <= "110001010010";
      when "00110001100" => color_data <= "110001010010";
      when "00110001101" => color_data <= "110001010010";
      when "00110001110" => color_data <= "110001010010";
      when "00110001111" => color_data <= "110001010010";
      when "00110010000" => color_data <= "110001010010";
      when "00110010001" => color_data <= "110001010010";
      when "00110010010" => color_data <= "110001010010";
      when "00110010011" => color_data <= "110001010010";
      when "00110010100" => color_data <= "110001010010";
      when "00110010101" => color_data <= "110101010010";
      when "00110010110" => color_data <= "101101000010";
      when "00110010111" => color_data <= "011000110010";
      when "00110011000" => color_data <= "101101000010";
      when "00110011001" => color_data <= "110101010010";
      when "00110011010" => color_data <= "110001010010";
      when "00110011011" => color_data <= "110001010010";
      when "00110011100" => color_data <= "110001010010";
      when "00110011101" => color_data <= "110001010010";
      when "00110011110" => color_data <= "110001010010";
      when "00110011111" => color_data <= "110001010010";
      when "00110100000" => color_data <= "110001010010";
      when "00110100001" => color_data <= "110001010010";
      when "00110100010" => color_data <= "110001010010";
      when "00110100011" => color_data <= "110001010010";
      when "00110100100" => color_data <= "110001010010";
      when "00110100101" => color_data <= "110001010010";
      when "00110100110" => color_data <= "110001010010";
      when "00110100111" => color_data <= "110001010010";
      when "00110101000" => color_data <= "110101010010";
      when "00110101001" => color_data <= "100001000010";
      when "00110101010" => color_data <= "011000110010";
      when "00110101011" => color_data <= "110101010010";
      when "00110101100" => color_data <= "110001010010";
      when "00110101101" => color_data <= "110001010010";
      when "00110101110" => color_data <= "110001010010";
      when "00110101111" => color_data <= "110001010010";
      when "00110110000" => color_data <= "110001010010";
      when "00110110001" => color_data <= "110001010010";
      when "00110110010" => color_data <= "110001010010";
      when "00110110011" => color_data <= "110001010010";
      when "00110110100" => color_data <= "110001010010";
      when "00110110101" => color_data <= "110001010010";
      when "00110110110" => color_data <= "110001010010";
      when "00110110111" => color_data <= "110001010010";
      when "00110111000" => color_data <= "110001010010";
      when "00110111001" => color_data <= "110001010010";
      when "00110111010" => color_data <= "110001010010";
      when "00110111011" => color_data <= "110101010010";
      when "00110111100" => color_data <= "011100110010";
      when "00110111101" => color_data <= "100101000010";
      when "00110111110" => color_data <= "110101010010";
      when "00110111111" => color_data <= "110001010010";
      when "00111000000" => color_data <= "100001000010";
      when "00111000001" => color_data <= "011100110010";
      when "00111000010" => color_data <= "100000110010";
      when "00111000011" => color_data <= "100000110010";
      when "00111000100" => color_data <= "011000110010";
      when "00111000101" => color_data <= "011100110010";
      when "00111000110" => color_data <= "100000110010";
      when "00111000111" => color_data <= "011100110010";
      when "00111001000" => color_data <= "011100110010";
      when "00111001001" => color_data <= "011100110010";
      when "00111001010" => color_data <= "011100110010";
      when "00111001011" => color_data <= "011100110010";
      when "00111001100" => color_data <= "011100110010";
      when "00111001101" => color_data <= "011100110010";
      when "00111001110" => color_data <= "011100110010";
      when "00111001111" => color_data <= "011100110010";
      when "00111010000" => color_data <= "011100110010";
      when "00111010001" => color_data <= "011100110010";
      when "00111010010" => color_data <= "011100110010";
      when "00111010011" => color_data <= "011100110010";
      when "00111010100" => color_data <= "011100110010";
      when "00111010101" => color_data <= "100000110010";
      when "00111010110" => color_data <= "011100110010";
      when "00111010111" => color_data <= "011000110010";
      when "00111011000" => color_data <= "011100110010";
      when "00111011001" => color_data <= "100000110010";
      when "00111011010" => color_data <= "011100110010";
      when "00111011011" => color_data <= "011100110010";
      when "00111011100" => color_data <= "011100110010";
      when "00111011101" => color_data <= "011100110010";
      when "00111011110" => color_data <= "011100110010";
      when "00111011111" => color_data <= "011100110010";
      when "00111100000" => color_data <= "011100110010";
      when "00111100001" => color_data <= "011100110010";
      when "00111100010" => color_data <= "011100110010";
      when "00111100011" => color_data <= "011100110010";
      when "00111100100" => color_data <= "011100110010";
      when "00111100101" => color_data <= "011100110010";
      when "00111100110" => color_data <= "011100110010";
      when "00111100111" => color_data <= "011100110010";
      when "00111101000" => color_data <= "100000110010";
      when "00111101001" => color_data <= "011000110010";
      when "00111101010" => color_data <= "011000110010";
      when "00111101011" => color_data <= "100000110010";
      when "00111101100" => color_data <= "100000110010";
      when "00111101101" => color_data <= "011100110010";
      when "00111101110" => color_data <= "011100110010";
      when "00111101111" => color_data <= "011100110010";
      when "00111110000" => color_data <= "011100110010";
      when "00111110001" => color_data <= "011100110010";
      when "00111110010" => color_data <= "011100110010";
      when "00111110011" => color_data <= "011100110010";
      when "00111110100" => color_data <= "011100110010";
      when "00111110101" => color_data <= "011100110010";
      when "00111110110" => color_data <= "011100110010";
      when "00111110111" => color_data <= "011100110010";
      when "00111111000" => color_data <= "011100110010";
      when "00111111001" => color_data <= "011100110010";
      when "00111111010" => color_data <= "011100110010";
      when "00111111011" => color_data <= "100000110010";
      when "00111111100" => color_data <= "011000110010";
      when "00111111101" => color_data <= "011100110010";
      when "00111111110" => color_data <= "100000110010";
      when "00111111111" => color_data <= "100001000010";
      when "01000000000" => color_data <= "101001010010";
      when "01000000001" => color_data <= "101001000010";
      when "01000000010" => color_data <= "101001000010";
      when "01000000011" => color_data <= "101001000010";
      when "01000000100" => color_data <= "101101000010";
      when "01000000101" => color_data <= "101101000010";
      when "01000000110" => color_data <= "101001000010";
      when "01000000111" => color_data <= "101001000010";
      when "01000001000" => color_data <= "101001000010";
      when "01000001001" => color_data <= "101001000010";
      when "01000001010" => color_data <= "101001000010";
      when "01000001011" => color_data <= "101001000010";
      when "01000001100" => color_data <= "101001000010";
      when "01000001101" => color_data <= "101001000010";
      when "01000001110" => color_data <= "010100110010";
      when "01000001111" => color_data <= "100101000010";
      when "01000010000" => color_data <= "101101000010";
      when "01000010001" => color_data <= "101001000010";
      when "01000010010" => color_data <= "101001000010";
      when "01000010011" => color_data <= "101001000010";
      when "01000010100" => color_data <= "101001000010";
      when "01000010101" => color_data <= "101001000010";
      when "01000010110" => color_data <= "101001000010";
      when "01000010111" => color_data <= "101101000010";
      when "01000011000" => color_data <= "101001000010";
      when "01000011001" => color_data <= "101001000010";
      when "01000011010" => color_data <= "101001000010";
      when "01000011011" => color_data <= "101001000010";
      when "01000011100" => color_data <= "101001000010";
      when "01000011101" => color_data <= "101001000010";
      when "01000011110" => color_data <= "101001000010";
      when "01000011111" => color_data <= "101101000010";
      when "01000100000" => color_data <= "100000110010";
      when "01000100001" => color_data <= "011000110010";
      when "01000100010" => color_data <= "101101000010";
      when "01000100011" => color_data <= "101001000010";
      when "01000100100" => color_data <= "101001000010";
      when "01000100101" => color_data <= "101001000010";
      when "01000100110" => color_data <= "101001000010";
      when "01000100111" => color_data <= "101001000010";
      when "01000101000" => color_data <= "101001000010";
      when "01000101001" => color_data <= "101101000010";
      when "01000101010" => color_data <= "101101000010";
      when "01000101011" => color_data <= "101001000010";
      when "01000101100" => color_data <= "101001000010";
      when "01000101101" => color_data <= "101001000010";
      when "01000101110" => color_data <= "101001000010";
      when "01000101111" => color_data <= "101001000010";
      when "01000110000" => color_data <= "101001000010";
      when "01000110001" => color_data <= "101001000010";
      when "01000110010" => color_data <= "101101000010";
      when "01000110011" => color_data <= "010100110010";
      when "01000110100" => color_data <= "011100110010";
      when "01000110101" => color_data <= "101101000010";
      when "01000110110" => color_data <= "101001000010";
      when "01000110111" => color_data <= "101001000010";
      when "01000111000" => color_data <= "101001000010";
      when "01000111001" => color_data <= "101001000010";
      when "01000111010" => color_data <= "101001000010";
      when "01000111011" => color_data <= "101001000010";
      when "01000111100" => color_data <= "101101000010";
      when "01000111101" => color_data <= "101101000010";
      when "01000111110" => color_data <= "101001000010";
      when "01000111111" => color_data <= "101001010010";
      when "01001000000" => color_data <= "110001010010";
      when "01001000001" => color_data <= "110001010010";
      when "01001000010" => color_data <= "110001010010";
      when "01001000011" => color_data <= "110001010010";
      when "01001000100" => color_data <= "110001010010";
      when "01001000101" => color_data <= "110001010010";
      when "01001000110" => color_data <= "110001010010";
      when "01001000111" => color_data <= "110001010010";
      when "01001001000" => color_data <= "110001010010";
      when "01001001001" => color_data <= "110001010010";
      when "01001001010" => color_data <= "110001010010";
      when "01001001011" => color_data <= "110001010010";
      when "01001001100" => color_data <= "110101010010";
      when "01001001101" => color_data <= "110001000010";
      when "01001001110" => color_data <= "011000110010";
      when "01001001111" => color_data <= "101101000010";
      when "01001010000" => color_data <= "110101010010";
      when "01001010001" => color_data <= "110001010010";
      when "01001010010" => color_data <= "110001010010";
      when "01001010011" => color_data <= "110001010010";
      when "01001010100" => color_data <= "110001010010";
      when "01001010101" => color_data <= "110001010010";
      when "01001010110" => color_data <= "110001010010";
      when "01001010111" => color_data <= "110001010010";
      when "01001011000" => color_data <= "110001010010";
      when "01001011001" => color_data <= "110001010010";
      when "01001011010" => color_data <= "110001010010";
      when "01001011011" => color_data <= "110001010010";
      when "01001011100" => color_data <= "110001010010";
      when "01001011101" => color_data <= "110001010010";
      when "01001011110" => color_data <= "110001010010";
      when "01001011111" => color_data <= "110101010010";
      when "01001100000" => color_data <= "100101000010";
      when "01001100001" => color_data <= "011100110010";
      when "01001100010" => color_data <= "110101010010";
      when "01001100011" => color_data <= "110001010010";
      when "01001100100" => color_data <= "110001010010";
      when "01001100101" => color_data <= "110001010010";
      when "01001100110" => color_data <= "110001010010";
      when "01001100111" => color_data <= "110001010010";
      when "01001101000" => color_data <= "110001010010";
      when "01001101001" => color_data <= "110001010010";
      when "01001101010" => color_data <= "110001010010";
      when "01001101011" => color_data <= "110001010010";
      when "01001101100" => color_data <= "110001010010";
      when "01001101101" => color_data <= "110001010010";
      when "01001101110" => color_data <= "110001010010";
      when "01001101111" => color_data <= "110001010010";
      when "01001110000" => color_data <= "110001010010";
      when "01001110001" => color_data <= "110001010010";
      when "01001110010" => color_data <= "110101010010";
      when "01001110011" => color_data <= "011000110010";
      when "01001110100" => color_data <= "100001000010";
      when "01001110101" => color_data <= "110101010010";
      when "01001110110" => color_data <= "110001010010";
      when "01001110111" => color_data <= "110001010010";
      when "01001111000" => color_data <= "110001010010";
      when "01001111001" => color_data <= "110001010010";
      when "01001111010" => color_data <= "110001010010";
      when "01001111011" => color_data <= "110001010010";
      when "01001111100" => color_data <= "110001010010";
      when "01001111101" => color_data <= "110001010010";
      when "01001111110" => color_data <= "110001010010";
      when "01001111111" => color_data <= "110001010010";
      when "01010000000" => color_data <= "110001010010";
      when "01010000001" => color_data <= "110001000010";
      when "01010000010" => color_data <= "110001000010";
      when "01010000011" => color_data <= "110001000010";
      when "01010000100" => color_data <= "110001000010";
      when "01010000101" => color_data <= "110001000010";
      when "01010000110" => color_data <= "110001000010";
      when "01010000111" => color_data <= "110001000010";
      when "01010001000" => color_data <= "110001000010";
      when "01010001001" => color_data <= "110001000010";
      when "01010001010" => color_data <= "110001000010";
      when "01010001011" => color_data <= "110001000010";
      when "01010001100" => color_data <= "110001010010";
      when "01010001101" => color_data <= "101101000010";
      when "01010001110" => color_data <= "011000110010";
      when "01010001111" => color_data <= "101001000010";
      when "01010010000" => color_data <= "110001010010";
      when "01010010001" => color_data <= "110001000010";
      when "01010010010" => color_data <= "110001000010";
      when "01010010011" => color_data <= "110001000010";
      when "01010010100" => color_data <= "110001000010";
      when "01010010101" => color_data <= "110001000010";
      when "01010010110" => color_data <= "110001000010";
      when "01010010111" => color_data <= "110001000010";
      when "01010011000" => color_data <= "110001000010";
      when "01010011001" => color_data <= "110001000010";
      when "01010011010" => color_data <= "110001000010";
      when "01010011011" => color_data <= "110001000010";
      when "01010011100" => color_data <= "110001000010";
      when "01010011101" => color_data <= "110001000010";
      when "01010011110" => color_data <= "110001000010";
      when "01010011111" => color_data <= "110101010010";
      when "01010100000" => color_data <= "100101000010";
      when "01010100001" => color_data <= "011100110010";
      when "01010100010" => color_data <= "110001010010";
      when "01010100011" => color_data <= "110001000010";
      when "01010100100" => color_data <= "110001000010";
      when "01010100101" => color_data <= "110001000010";
      when "01010100110" => color_data <= "110001000010";
      when "01010100111" => color_data <= "110001000010";
      when "01010101000" => color_data <= "110001000010";
      when "01010101001" => color_data <= "110001000010";
      when "01010101010" => color_data <= "110001000010";
      when "01010101011" => color_data <= "110001000010";
      when "01010101100" => color_data <= "110001000010";
      when "01010101101" => color_data <= "110001000010";
      when "01010101110" => color_data <= "110001000010";
      when "01010101111" => color_data <= "110001000010";
      when "01010110000" => color_data <= "110001000010";
      when "01010110001" => color_data <= "110001000010";
      when "01010110010" => color_data <= "110001010010";
      when "01010110011" => color_data <= "011000110010";
      when "01010110100" => color_data <= "100001000010";
      when "01010110101" => color_data <= "110101010010";
      when "01010110110" => color_data <= "110001000010";
      when "01010110111" => color_data <= "110001000010";
      when "01010111000" => color_data <= "110001000010";
      when "01010111001" => color_data <= "110001000010";
      when "01010111010" => color_data <= "110001000010";
      when "01010111011" => color_data <= "110001000010";
      when "01010111100" => color_data <= "110001000010";
      when "01010111101" => color_data <= "110001000010";
      when "01010111110" => color_data <= "110001000010";
      when "01010111111" => color_data <= "110001010010";
      when "01011000000" => color_data <= "110001010010";
      when "01011000001" => color_data <= "110001000010";
      when "01011000010" => color_data <= "110001000010";
      when "01011000011" => color_data <= "110001000010";
      when "01011000100" => color_data <= "110001000010";
      when "01011000101" => color_data <= "110001000010";
      when "01011000110" => color_data <= "110001000010";
      when "01011000111" => color_data <= "110001000010";
      when "01011001000" => color_data <= "110001000010";
      when "01011001001" => color_data <= "110001000010";
      when "01011001010" => color_data <= "110001000010";
      when "01011001011" => color_data <= "110001000010";
      when "01011001100" => color_data <= "110001010010";
      when "01011001101" => color_data <= "101101000010";
      when "01011001110" => color_data <= "011000110010";
      when "01011001111" => color_data <= "101001000010";
      when "01011010000" => color_data <= "110001010010";
      when "01011010001" => color_data <= "110001000010";
      when "01011010010" => color_data <= "110001000010";
      when "01011010011" => color_data <= "110001000010";
      when "01011010100" => color_data <= "110001000010";
      when "01011010101" => color_data <= "110001000010";
      when "01011010110" => color_data <= "110001000010";
      when "01011010111" => color_data <= "110001000010";
      when "01011011000" => color_data <= "110001000010";
      when "01011011001" => color_data <= "110001000010";
      when "01011011010" => color_data <= "110001000010";
      when "01011011011" => color_data <= "110001000010";
      when "01011011100" => color_data <= "110001000010";
      when "01011011101" => color_data <= "110001000010";
      when "01011011110" => color_data <= "110001000010";
      when "01011011111" => color_data <= "110101010010";
      when "01011100000" => color_data <= "100101000010";
      when "01011100001" => color_data <= "011100110010";
      when "01011100010" => color_data <= "110001010010";
      when "01011100011" => color_data <= "110001000010";
      when "01011100100" => color_data <= "110001000010";
      when "01011100101" => color_data <= "110001000010";
      when "01011100110" => color_data <= "110001000010";
      when "01011100111" => color_data <= "110001000010";
      when "01011101000" => color_data <= "110001000010";
      when "01011101001" => color_data <= "110001000010";
      when "01011101010" => color_data <= "110001000010";
      when "01011101011" => color_data <= "110001000010";
      when "01011101100" => color_data <= "110001000010";
      when "01011101101" => color_data <= "110001000010";
      when "01011101110" => color_data <= "110001000010";
      when "01011101111" => color_data <= "110001000010";
      when "01011110000" => color_data <= "110001000010";
      when "01011110001" => color_data <= "110001000010";
      when "01011110010" => color_data <= "110001010010";
      when "01011110011" => color_data <= "011000110010";
      when "01011110100" => color_data <= "100001000010";
      when "01011110101" => color_data <= "110101010010";
      when "01011110110" => color_data <= "110001000010";
      when "01011110111" => color_data <= "110001000010";
      when "01011111000" => color_data <= "110001000010";
      when "01011111001" => color_data <= "110001000010";
      when "01011111010" => color_data <= "110001000010";
      when "01011111011" => color_data <= "110001000010";
      when "01011111100" => color_data <= "110001000010";
      when "01011111101" => color_data <= "110001000010";
      when "01011111110" => color_data <= "110001000010";
      when "01011111111" => color_data <= "110001010010";
      when "01100000000" => color_data <= "110001010010";
      when "01100000001" => color_data <= "110001000010";
      when "01100000010" => color_data <= "110001000010";
      when "01100000011" => color_data <= "110001000010";
      when "01100000100" => color_data <= "110001000010";
      when "01100000101" => color_data <= "110001000010";
      when "01100000110" => color_data <= "110001000010";
      when "01100000111" => color_data <= "110001000010";
      when "01100001000" => color_data <= "110001000010";
      when "01100001001" => color_data <= "110001000010";
      when "01100001010" => color_data <= "110001000010";
      when "01100001011" => color_data <= "110001000010";
      when "01100001100" => color_data <= "110001010010";
      when "01100001101" => color_data <= "101101000010";
      when "01100001110" => color_data <= "011000110010";
      when "01100001111" => color_data <= "101001000010";
      when "01100010000" => color_data <= "110001010010";
      when "01100010001" => color_data <= "110001000010";
      when "01100010010" => color_data <= "110001000010";
      when "01100010011" => color_data <= "110001000010";
      when "01100010100" => color_data <= "110001000010";
      when "01100010101" => color_data <= "110001000010";
      when "01100010110" => color_data <= "110001000010";
      when "01100010111" => color_data <= "110001000010";
      when "01100011000" => color_data <= "110001000010";
      when "01100011001" => color_data <= "110001000010";
      when "01100011010" => color_data <= "110001000010";
      when "01100011011" => color_data <= "110001000010";
      when "01100011100" => color_data <= "110001000010";
      when "01100011101" => color_data <= "110001000010";
      when "01100011110" => color_data <= "110001000010";
      when "01100011111" => color_data <= "110101010010";
      when "01100100000" => color_data <= "100101000010";
      when "01100100001" => color_data <= "011100110010";
      when "01100100010" => color_data <= "110001010010";
      when "01100100011" => color_data <= "110001000010";
      when "01100100100" => color_data <= "110001000010";
      when "01100100101" => color_data <= "110001000010";
      when "01100100110" => color_data <= "110001000010";
      when "01100100111" => color_data <= "110001000010";
      when "01100101000" => color_data <= "110001000010";
      when "01100101001" => color_data <= "110001000010";
      when "01100101010" => color_data <= "110001000010";
      when "01100101011" => color_data <= "110001000010";
      when "01100101100" => color_data <= "110001000010";
      when "01100101101" => color_data <= "110001000010";
      when "01100101110" => color_data <= "110001000010";
      when "01100101111" => color_data <= "110001000010";
      when "01100110000" => color_data <= "110001000010";
      when "01100110001" => color_data <= "110001000010";
      when "01100110010" => color_data <= "110001010010";
      when "01100110011" => color_data <= "011000110010";
      when "01100110100" => color_data <= "100001000010";
      when "01100110101" => color_data <= "110101010010";
      when "01100110110" => color_data <= "110001000010";
      when "01100110111" => color_data <= "110001000010";
      when "01100111000" => color_data <= "110001000010";
      when "01100111001" => color_data <= "110001000010";
      when "01100111010" => color_data <= "110001000010";
      when "01100111011" => color_data <= "110001000010";
      when "01100111100" => color_data <= "110001000010";
      when "01100111101" => color_data <= "110001000010";
      when "01100111110" => color_data <= "110001000010";
      when "01100111111" => color_data <= "110001010010";
      when "01101000000" => color_data <= "110001010010";
      when "01101000001" => color_data <= "110001000010";
      when "01101000010" => color_data <= "110001000010";
      when "01101000011" => color_data <= "110001000010";
      when "01101000100" => color_data <= "110001000010";
      when "01101000101" => color_data <= "110001000010";
      when "01101000110" => color_data <= "110001000010";
      when "01101000111" => color_data <= "110001000010";
      when "01101001000" => color_data <= "110001000010";
      when "01101001001" => color_data <= "110001000010";
      when "01101001010" => color_data <= "110001000010";
      when "01101001011" => color_data <= "110001000010";
      when "01101001100" => color_data <= "110001010010";
      when "01101001101" => color_data <= "101101000010";
      when "01101001110" => color_data <= "011000110010";
      when "01101001111" => color_data <= "101001000010";
      when "01101010000" => color_data <= "110001010010";
      when "01101010001" => color_data <= "110001000010";
      when "01101010010" => color_data <= "110001000010";
      when "01101010011" => color_data <= "110001000010";
      when "01101010100" => color_data <= "110001000010";
      when "01101010101" => color_data <= "110001000010";
      when "01101010110" => color_data <= "110001000010";
      when "01101010111" => color_data <= "110001000010";
      when "01101011000" => color_data <= "110001000010";
      when "01101011001" => color_data <= "110001000010";
      when "01101011010" => color_data <= "110001000010";
      when "01101011011" => color_data <= "110001000010";
      when "01101011100" => color_data <= "110001000010";
      when "01101011101" => color_data <= "110001000010";
      when "01101011110" => color_data <= "110001000010";
      when "01101011111" => color_data <= "110101010010";
      when "01101100000" => color_data <= "100101000010";
      when "01101100001" => color_data <= "011100110010";
      when "01101100010" => color_data <= "110001010010";
      when "01101100011" => color_data <= "110001000010";
      when "01101100100" => color_data <= "110001000010";
      when "01101100101" => color_data <= "110001000010";
      when "01101100110" => color_data <= "110001000010";
      when "01101100111" => color_data <= "110001000010";
      when "01101101000" => color_data <= "110001000010";
      when "01101101001" => color_data <= "110001000010";
      when "01101101010" => color_data <= "110001000010";
      when "01101101011" => color_data <= "110001000010";
      when "01101101100" => color_data <= "110001000010";
      when "01101101101" => color_data <= "110001000010";
      when "01101101110" => color_data <= "110001000010";
      when "01101101111" => color_data <= "110001000010";
      when "01101110000" => color_data <= "110001000010";
      when "01101110001" => color_data <= "110001000010";
      when "01101110010" => color_data <= "110001010010";
      when "01101110011" => color_data <= "011000110010";
      when "01101110100" => color_data <= "100001000010";
      when "01101110101" => color_data <= "110101010010";
      when "01101110110" => color_data <= "110001000010";
      when "01101110111" => color_data <= "110001000010";
      when "01101111000" => color_data <= "110001000010";
      when "01101111001" => color_data <= "110001000010";
      when "01101111010" => color_data <= "110001000010";
      when "01101111011" => color_data <= "110001000010";
      when "01101111100" => color_data <= "110001000010";
      when "01101111101" => color_data <= "110001000010";
      when "01101111110" => color_data <= "110001000010";
      when "01101111111" => color_data <= "110001010010";
      when "01110000000" => color_data <= "110101010010";
      when "01110000001" => color_data <= "110101010010";
      when "01110000010" => color_data <= "110101010010";
      when "01110000011" => color_data <= "110101010010";
      when "01110000100" => color_data <= "110101010010";
      when "01110000101" => color_data <= "110101010010";
      when "01110000110" => color_data <= "110101010010";
      when "01110000111" => color_data <= "110101010010";
      when "01110001000" => color_data <= "110101010010";
      when "01110001001" => color_data <= "110101010010";
      when "01110001010" => color_data <= "110101010010";
      when "01110001011" => color_data <= "110101010010";
      when "01110001100" => color_data <= "110101010010";
      when "01110001101" => color_data <= "110001010010";
      when "01110001110" => color_data <= "011000110010";
      when "01110001111" => color_data <= "101101000010";
      when "01110010000" => color_data <= "110101010010";
      when "01110010001" => color_data <= "110101010010";
      when "01110010010" => color_data <= "110101010010";
      when "01110010011" => color_data <= "110101010010";
      when "01110010100" => color_data <= "110101010010";
      when "01110010101" => color_data <= "110101010010";
      when "01110010110" => color_data <= "110101010010";
      when "01110010111" => color_data <= "110101010010";
      when "01110011000" => color_data <= "110101010010";
      when "01110011001" => color_data <= "110101010010";
      when "01110011010" => color_data <= "110101010010";
      when "01110011011" => color_data <= "110101010010";
      when "01110011100" => color_data <= "110101010010";
      when "01110011101" => color_data <= "110101010010";
      when "01110011110" => color_data <= "110101010010";
      when "01110011111" => color_data <= "111001010010";
      when "01110100000" => color_data <= "100101000010";
      when "01110100001" => color_data <= "011100110010";
      when "01110100010" => color_data <= "111001010010";
      when "01110100011" => color_data <= "110101010010";
      when "01110100100" => color_data <= "110101010010";
      when "01110100101" => color_data <= "110101010010";
      when "01110100110" => color_data <= "110101010010";
      when "01110100111" => color_data <= "110101010010";
      when "01110101000" => color_data <= "110101010010";
      when "01110101001" => color_data <= "110101010010";
      when "01110101010" => color_data <= "110101010010";
      when "01110101011" => color_data <= "110101010010";
      when "01110101100" => color_data <= "110101010010";
      when "01110101101" => color_data <= "110101010010";
      when "01110101110" => color_data <= "110101010010";
      when "01110101111" => color_data <= "110101010010";
      when "01110110000" => color_data <= "110101010010";
      when "01110110001" => color_data <= "110101010010";
      when "01110110010" => color_data <= "110101010010";
      when "01110110011" => color_data <= "011000110010";
      when "01110110100" => color_data <= "100001000010";
      when "01110110101" => color_data <= "111001010010";
      when "01110110110" => color_data <= "110101010010";
      when "01110110111" => color_data <= "110101010010";
      when "01110111000" => color_data <= "110101010010";
      when "01110111001" => color_data <= "110101010010";
      when "01110111010" => color_data <= "110101010010";
      when "01110111011" => color_data <= "110101010010";
      when "01110111100" => color_data <= "110101010010";
      when "01110111101" => color_data <= "110101010010";
      when "01110111110" => color_data <= "110101010010";
      when "01110111111" => color_data <= "110101010010";
      when "01111000000" => color_data <= "100101000010";
      when "01111000001" => color_data <= "100001000010";
      when "01111000010" => color_data <= "100001000010";
      when "01111000011" => color_data <= "100001000010";
      when "01111000100" => color_data <= "100001000010";
      when "01111000101" => color_data <= "100001000010";
      when "01111000110" => color_data <= "100001000010";
      when "01111000111" => color_data <= "100001000010";
      when "01111001000" => color_data <= "100101000010";
      when "01111001001" => color_data <= "100101000010";
      when "01111001010" => color_data <= "100001000010";
      when "01111001011" => color_data <= "100001000010";
      when "01111001100" => color_data <= "100101000010";
      when "01111001101" => color_data <= "100001000010";
      when "01111001110" => color_data <= "010100110010";
      when "01111001111" => color_data <= "100000110010";
      when "01111010000" => color_data <= "100101000010";
      when "01111010001" => color_data <= "100001000010";
      when "01111010010" => color_data <= "100001000010";
      when "01111010011" => color_data <= "100001000010";
      when "01111010100" => color_data <= "100001000010";
      when "01111010101" => color_data <= "100001000010";
      when "01111010110" => color_data <= "100001000010";
      when "01111010111" => color_data <= "100001000010";
      when "01111011000" => color_data <= "100001000010";
      when "01111011001" => color_data <= "100001000010";
      when "01111011010" => color_data <= "100001000010";
      when "01111011011" => color_data <= "100101000010";
      when "01111011100" => color_data <= "100101000010";
      when "01111011101" => color_data <= "100001000010";
      when "01111011110" => color_data <= "100001000010";
      when "01111011111" => color_data <= "100101000010";
      when "01111100000" => color_data <= "011100110010";
      when "01111100001" => color_data <= "011000110010";
      when "01111100010" => color_data <= "100101000010";
      when "01111100011" => color_data <= "100001000010";
      when "01111100100" => color_data <= "100001000010";
      when "01111100101" => color_data <= "100001000010";
      when "01111100110" => color_data <= "100001000010";
      when "01111100111" => color_data <= "100001000010";
      when "01111101000" => color_data <= "100001000010";
      when "01111101001" => color_data <= "100001000010";
      when "01111101010" => color_data <= "100001000010";
      when "01111101011" => color_data <= "100001000010";
      when "01111101100" => color_data <= "100001000010";
      when "01111101101" => color_data <= "100101000010";
      when "01111101110" => color_data <= "100101000010";
      when "01111101111" => color_data <= "100001000010";
      when "01111110000" => color_data <= "100001000010";
      when "01111110001" => color_data <= "100001000010";
      when "01111110010" => color_data <= "100101000010";
      when "01111110011" => color_data <= "010100110010";
      when "01111110100" => color_data <= "011000110010";
      when "01111110101" => color_data <= "100101000010";
      when "01111110110" => color_data <= "100001000010";
      when "01111110111" => color_data <= "100001000010";
      when "01111111000" => color_data <= "100001000010";
      when "01111111001" => color_data <= "100001000010";
      when "01111111010" => color_data <= "100001000010";
      when "01111111011" => color_data <= "100001000010";
      when "01111111100" => color_data <= "100001000010";
      when "01111111101" => color_data <= "100001000010";
      when "01111111110" => color_data <= "100001000010";
      when "01111111111" => color_data <= "100101000010";
      when "10000000000" => color_data <= "100101000010";
      when "10000000001" => color_data <= "100101000010";
      when "10000000010" => color_data <= "100101000010";
      when "10000000011" => color_data <= "100101000010";
      when "10000000100" => color_data <= "100101000010";
      when "10000000101" => color_data <= "100101000010";
      when "10000000110" => color_data <= "100101000010";
      when "10000000111" => color_data <= "101001000010";
      when "10000001000" => color_data <= "011000110010";
      when "10000001001" => color_data <= "011000110010";
      when "10000001010" => color_data <= "100101000010";
      when "10000001011" => color_data <= "100101000010";
      when "10000001100" => color_data <= "100101000010";
      when "10000001101" => color_data <= "100101000010";
      when "10000001110" => color_data <= "101001000010";
      when "10000001111" => color_data <= "100101000010";
      when "10000010000" => color_data <= "100101000010";
      when "10000010001" => color_data <= "100101000010";
      when "10000010010" => color_data <= "100101000010";
      when "10000010011" => color_data <= "100101000010";
      when "10000010100" => color_data <= "100101000010";
      when "10000010101" => color_data <= "100101000010";
      when "10000010110" => color_data <= "100101000010";
      when "10000010111" => color_data <= "100101000010";
      when "10000011000" => color_data <= "100101000010";
      when "10000011001" => color_data <= "100101000010";
      when "10000011010" => color_data <= "100101000010";
      when "10000011011" => color_data <= "010100110010";
      when "10000011100" => color_data <= "011100110010";
      when "10000011101" => color_data <= "100101000010";
      when "10000011110" => color_data <= "100101000010";
      when "10000011111" => color_data <= "100101000010";
      when "10000100000" => color_data <= "100101000010";
      when "10000100001" => color_data <= "101001000010";
      when "10000100010" => color_data <= "100101000010";
      when "10000100011" => color_data <= "100101000010";
      when "10000100100" => color_data <= "100101000010";
      when "10000100101" => color_data <= "100101000010";
      when "10000100110" => color_data <= "100101000010";
      when "10000100111" => color_data <= "100101000010";
      when "10000101000" => color_data <= "100101000010";
      when "10000101001" => color_data <= "100101000010";
      when "10000101010" => color_data <= "100101000010";
      when "10000101011" => color_data <= "100101000010";
      when "10000101100" => color_data <= "100101000010";
      when "10000101101" => color_data <= "100000110010";
      when "10000101110" => color_data <= "010100110010";
      when "10000101111" => color_data <= "100101000010";
      when "10000110000" => color_data <= "100101000010";
      when "10000110001" => color_data <= "100101000010";
      when "10000110010" => color_data <= "100101000010";
      when "10000110011" => color_data <= "101001000010";
      when "10000110100" => color_data <= "100101000010";
      when "10000110101" => color_data <= "100101000010";
      when "10000110110" => color_data <= "100101000010";
      when "10000110111" => color_data <= "100101000010";
      when "10000111000" => color_data <= "100101000010";
      when "10000111001" => color_data <= "100101000010";
      when "10000111010" => color_data <= "100101000010";
      when "10000111011" => color_data <= "100101000010";
      when "10000111100" => color_data <= "100101000010";
      when "10000111101" => color_data <= "100101000010";
      when "10000111110" => color_data <= "100101000010";
      when "10000111111" => color_data <= "100101000010";
      when "10001000000" => color_data <= "110101010010";
      when "10001000001" => color_data <= "110101010010";
      when "10001000010" => color_data <= "110101010010";
      when "10001000011" => color_data <= "110101010010";
      when "10001000100" => color_data <= "110101010010";
      when "10001000101" => color_data <= "110101010010";
      when "10001000110" => color_data <= "110101010010";
      when "10001000111" => color_data <= "111001010010";
      when "10001001000" => color_data <= "100001000010";
      when "10001001001" => color_data <= "011100110010";
      when "10001001010" => color_data <= "111001010010";
      when "10001001011" => color_data <= "110101010010";
      when "10001001100" => color_data <= "110101010010";
      when "10001001101" => color_data <= "110101010010";
      when "10001001110" => color_data <= "110101010010";
      when "10001001111" => color_data <= "110101010010";
      when "10001010000" => color_data <= "110101010010";
      when "10001010001" => color_data <= "110101010010";
      when "10001010010" => color_data <= "110101010010";
      when "10001010011" => color_data <= "110101010010";
      when "10001010100" => color_data <= "110101010010";
      when "10001010101" => color_data <= "110101010010";
      when "10001010110" => color_data <= "110101010010";
      when "10001010111" => color_data <= "110101010010";
      when "10001011000" => color_data <= "110101010010";
      when "10001011001" => color_data <= "110101010010";
      when "10001011010" => color_data <= "110101010010";
      when "10001011011" => color_data <= "011100110010";
      when "10001011100" => color_data <= "101001000010";
      when "10001011101" => color_data <= "111001010010";
      when "10001011110" => color_data <= "110101010010";
      when "10001011111" => color_data <= "110101010010";
      when "10001100000" => color_data <= "110101010010";
      when "10001100001" => color_data <= "110101010010";
      when "10001100010" => color_data <= "110101010010";
      when "10001100011" => color_data <= "110101010010";
      when "10001100100" => color_data <= "110101010010";
      when "10001100101" => color_data <= "110101010010";
      when "10001100110" => color_data <= "110101010010";
      when "10001100111" => color_data <= "110101010010";
      when "10001101000" => color_data <= "110101010010";
      when "10001101001" => color_data <= "110101010010";
      when "10001101010" => color_data <= "110101010010";
      when "10001101011" => color_data <= "110101010010";
      when "10001101100" => color_data <= "111001010010";
      when "10001101101" => color_data <= "101001000010";
      when "10001101110" => color_data <= "011000110010";
      when "10001101111" => color_data <= "110101010010";
      when "10001110000" => color_data <= "110101010010";
      when "10001110001" => color_data <= "110101010010";
      when "10001110010" => color_data <= "110101010010";
      when "10001110011" => color_data <= "110101010010";
      when "10001110100" => color_data <= "110101010010";
      when "10001110101" => color_data <= "110101010010";
      when "10001110110" => color_data <= "110101010010";
      when "10001110111" => color_data <= "110101010010";
      when "10001111000" => color_data <= "110101010010";
      when "10001111001" => color_data <= "110101010010";
      when "10001111010" => color_data <= "110101010010";
      when "10001111011" => color_data <= "110101010010";
      when "10001111100" => color_data <= "110101010010";
      when "10001111101" => color_data <= "110101010010";
      when "10001111110" => color_data <= "110101010010";
      when "10001111111" => color_data <= "110101010010";
      when "10010000000" => color_data <= "110001010010";
      when "10010000001" => color_data <= "110001000010";
      when "10010000010" => color_data <= "110001000010";
      when "10010000011" => color_data <= "110001000010";
      when "10010000100" => color_data <= "110001000010";
      when "10010000101" => color_data <= "110001000010";
      when "10010000110" => color_data <= "110001000010";
      when "10010000111" => color_data <= "110101010010";
      when "10010001000" => color_data <= "100001000010";
      when "10010001001" => color_data <= "011100110010";
      when "10010001010" => color_data <= "110101010010";
      when "10010001011" => color_data <= "110001000010";
      when "10010001100" => color_data <= "110001000010";
      when "10010001101" => color_data <= "110001000010";
      when "10010001110" => color_data <= "110001000010";
      when "10010001111" => color_data <= "110001000010";
      when "10010010000" => color_data <= "110001000010";
      when "10010010001" => color_data <= "110001000010";
      when "10010010010" => color_data <= "110001000010";
      when "10010010011" => color_data <= "110001000010";
      when "10010010100" => color_data <= "110001000010";
      when "10010010101" => color_data <= "110001000010";
      when "10010010110" => color_data <= "110001000010";
      when "10010010111" => color_data <= "110001000010";
      when "10010011000" => color_data <= "110001000010";
      when "10010011001" => color_data <= "110001000010";
      when "10010011010" => color_data <= "110001010010";
      when "10010011011" => color_data <= "011100110010";
      when "10010011100" => color_data <= "100101000010";
      when "10010011101" => color_data <= "110101010010";
      when "10010011110" => color_data <= "110001000010";
      when "10010011111" => color_data <= "110001000010";
      when "10010100000" => color_data <= "110001000010";
      when "10010100001" => color_data <= "110001000010";
      when "10010100010" => color_data <= "110001000010";
      when "10010100011" => color_data <= "110001000010";
      when "10010100100" => color_data <= "110001000010";
      when "10010100101" => color_data <= "110001000010";
      when "10010100110" => color_data <= "110001000010";
      when "10010100111" => color_data <= "110001000010";
      when "10010101000" => color_data <= "110001000010";
      when "10010101001" => color_data <= "110001000010";
      when "10010101010" => color_data <= "110001000010";
      when "10010101011" => color_data <= "110001000010";
      when "10010101100" => color_data <= "110101010010";
      when "10010101101" => color_data <= "101001000010";
      when "10010101110" => color_data <= "011000110010";
      when "10010101111" => color_data <= "110001000010";
      when "10010110000" => color_data <= "110001010010";
      when "10010110001" => color_data <= "110001000010";
      when "10010110010" => color_data <= "110001000010";
      when "10010110011" => color_data <= "110001000010";
      when "10010110100" => color_data <= "110001000010";
      when "10010110101" => color_data <= "110001000010";
      when "10010110110" => color_data <= "110001000010";
      when "10010110111" => color_data <= "110001000010";
      when "10010111000" => color_data <= "110001000010";
      when "10010111001" => color_data <= "110001000010";
      when "10010111010" => color_data <= "110001000010";
      when "10010111011" => color_data <= "110001000010";
      when "10010111100" => color_data <= "110001000010";
      when "10010111101" => color_data <= "110001000010";
      when "10010111110" => color_data <= "110001000010";
      when "10010111111" => color_data <= "110001010010";
      when "10011000000" => color_data <= "110001010010";
      when "10011000001" => color_data <= "110001000010";
      when "10011000010" => color_data <= "110001000010";
      when "10011000011" => color_data <= "110001000010";
      when "10011000100" => color_data <= "110001000010";
      when "10011000101" => color_data <= "110001000010";
      when "10011000110" => color_data <= "110001000010";
      when "10011000111" => color_data <= "110101010010";
      when "10011001000" => color_data <= "100001000010";
      when "10011001001" => color_data <= "011100110010";
      when "10011001010" => color_data <= "110101010010";
      when "10011001011" => color_data <= "110001000010";
      when "10011001100" => color_data <= "110001000010";
      when "10011001101" => color_data <= "110001000010";
      when "10011001110" => color_data <= "110001000010";
      when "10011001111" => color_data <= "110001000010";
      when "10011010000" => color_data <= "110001000010";
      when "10011010001" => color_data <= "110001000010";
      when "10011010010" => color_data <= "110001000010";
      when "10011010011" => color_data <= "110001000010";
      when "10011010100" => color_data <= "110001000010";
      when "10011010101" => color_data <= "110001000010";
      when "10011010110" => color_data <= "110001000010";
      when "10011010111" => color_data <= "110001000010";
      when "10011011000" => color_data <= "110001000010";
      when "10011011001" => color_data <= "110001000010";
      when "10011011010" => color_data <= "110001010010";
      when "10011011011" => color_data <= "011100110010";
      when "10011011100" => color_data <= "100101000010";
      when "10011011101" => color_data <= "110101010010";
      when "10011011110" => color_data <= "110001000010";
      when "10011011111" => color_data <= "110001000010";
      when "10011100000" => color_data <= "110001000010";
      when "10011100001" => color_data <= "110001000010";
      when "10011100010" => color_data <= "110001000010";
      when "10011100011" => color_data <= "110001000010";
      when "10011100100" => color_data <= "110001000010";
      when "10011100101" => color_data <= "110001000010";
      when "10011100110" => color_data <= "110001000010";
      when "10011100111" => color_data <= "110001000010";
      when "10011101000" => color_data <= "110001000010";
      when "10011101001" => color_data <= "110001000010";
      when "10011101010" => color_data <= "110001000010";
      when "10011101011" => color_data <= "110001000010";
      when "10011101100" => color_data <= "110101010010";
      when "10011101101" => color_data <= "101001000010";
      when "10011101110" => color_data <= "011000110010";
      when "10011101111" => color_data <= "110001000010";
      when "10011110000" => color_data <= "110001010010";
      when "10011110001" => color_data <= "110001000010";
      when "10011110010" => color_data <= "110001000010";
      when "10011110011" => color_data <= "110001000010";
      when "10011110100" => color_data <= "110001000010";
      when "10011110101" => color_data <= "110001000010";
      when "10011110110" => color_data <= "110001000010";
      when "10011110111" => color_data <= "110001000010";
      when "10011111000" => color_data <= "110001000010";
      when "10011111001" => color_data <= "110001000010";
      when "10011111010" => color_data <= "110001000010";
      when "10011111011" => color_data <= "110001000010";
      when "10011111100" => color_data <= "110001000010";
      when "10011111101" => color_data <= "110001000010";
      when "10011111110" => color_data <= "110001000010";
      when "10011111111" => color_data <= "110001010010";
      when "10100000000" => color_data <= "110001010010";
      when "10100000001" => color_data <= "110001000010";
      when "10100000010" => color_data <= "110001000010";
      when "10100000011" => color_data <= "110001000010";
      when "10100000100" => color_data <= "110001000010";
      when "10100000101" => color_data <= "110001000010";
      when "10100000110" => color_data <= "110001000010";
      when "10100000111" => color_data <= "110101010010";
      when "10100001000" => color_data <= "100001000010";
      when "10100001001" => color_data <= "011100110010";
      when "10100001010" => color_data <= "110101010010";
      when "10100001011" => color_data <= "110001000010";
      when "10100001100" => color_data <= "110001000010";
      when "10100001101" => color_data <= "110001000010";
      when "10100001110" => color_data <= "110001000010";
      when "10100001111" => color_data <= "110001000010";
      when "10100010000" => color_data <= "110001000010";
      when "10100010001" => color_data <= "110001000010";
      when "10100010010" => color_data <= "110001000010";
      when "10100010011" => color_data <= "110001000010";
      when "10100010100" => color_data <= "110001000010";
      when "10100010101" => color_data <= "110001000010";
      when "10100010110" => color_data <= "110001000010";
      when "10100010111" => color_data <= "110001000010";
      when "10100011000" => color_data <= "110001000010";
      when "10100011001" => color_data <= "110001000010";
      when "10100011010" => color_data <= "110001010010";
      when "10100011011" => color_data <= "011100110010";
      when "10100011100" => color_data <= "100101000010";
      when "10100011101" => color_data <= "110101010010";
      when "10100011110" => color_data <= "110001000010";
      when "10100011111" => color_data <= "110001000010";
      when "10100100000" => color_data <= "110001000010";
      when "10100100001" => color_data <= "110001000010";
      when "10100100010" => color_data <= "110001000010";
      when "10100100011" => color_data <= "110001000010";
      when "10100100100" => color_data <= "110001000010";
      when "10100100101" => color_data <= "110001000010";
      when "10100100110" => color_data <= "110001000010";
      when "10100100111" => color_data <= "110001000010";
      when "10100101000" => color_data <= "110001000010";
      when "10100101001" => color_data <= "110001000010";
      when "10100101010" => color_data <= "110001000010";
      when "10100101011" => color_data <= "110001000010";
      when "10100101100" => color_data <= "110101010010";
      when "10100101101" => color_data <= "101001000010";
      when "10100101110" => color_data <= "011000110010";
      when "10100101111" => color_data <= "110001000010";
      when "10100110000" => color_data <= "110001010010";
      when "10100110001" => color_data <= "110001000010";
      when "10100110010" => color_data <= "110001000010";
      when "10100110011" => color_data <= "110001000010";
      when "10100110100" => color_data <= "110001000010";
      when "10100110101" => color_data <= "110001000010";
      when "10100110110" => color_data <= "110001000010";
      when "10100110111" => color_data <= "110001000010";
      when "10100111000" => color_data <= "110001000010";
      when "10100111001" => color_data <= "110001000010";
      when "10100111010" => color_data <= "110001000010";
      when "10100111011" => color_data <= "110001000010";
      when "10100111100" => color_data <= "110001000010";
      when "10100111101" => color_data <= "110001000010";
      when "10100111110" => color_data <= "110001000010";
      when "10100111111" => color_data <= "110001010010";
      when "10101000000" => color_data <= "110001010010";
      when "10101000001" => color_data <= "110001000010";
      when "10101000010" => color_data <= "110001000010";
      when "10101000011" => color_data <= "110001000010";
      when "10101000100" => color_data <= "110001000010";
      when "10101000101" => color_data <= "110001000010";
      when "10101000110" => color_data <= "110001000010";
      when "10101000111" => color_data <= "110101010010";
      when "10101001000" => color_data <= "100001000010";
      when "10101001001" => color_data <= "011100110010";
      when "10101001010" => color_data <= "110101010010";
      when "10101001011" => color_data <= "110001000010";
      when "10101001100" => color_data <= "110001000010";
      when "10101001101" => color_data <= "110001000010";
      when "10101001110" => color_data <= "110001000010";
      when "10101001111" => color_data <= "110001000010";
      when "10101010000" => color_data <= "110001000010";
      when "10101010001" => color_data <= "110001000010";
      when "10101010010" => color_data <= "110001000010";
      when "10101010011" => color_data <= "110001000010";
      when "10101010100" => color_data <= "110001000010";
      when "10101010101" => color_data <= "110001000010";
      when "10101010110" => color_data <= "110001000010";
      when "10101010111" => color_data <= "110001000010";
      when "10101011000" => color_data <= "110001000010";
      when "10101011001" => color_data <= "110001000010";
      when "10101011010" => color_data <= "110001010010";
      when "10101011011" => color_data <= "011100110010";
      when "10101011100" => color_data <= "100101000010";
      when "10101011101" => color_data <= "110101010010";
      when "10101011110" => color_data <= "110001000010";
      when "10101011111" => color_data <= "110001000010";
      when "10101100000" => color_data <= "110001000010";
      when "10101100001" => color_data <= "110001000010";
      when "10101100010" => color_data <= "110001000010";
      when "10101100011" => color_data <= "110001000010";
      when "10101100100" => color_data <= "110001000010";
      when "10101100101" => color_data <= "110001000010";
      when "10101100110" => color_data <= "110001000010";
      when "10101100111" => color_data <= "110001000010";
      when "10101101000" => color_data <= "110001000010";
      when "10101101001" => color_data <= "110001000010";
      when "10101101010" => color_data <= "110001000010";
      when "10101101011" => color_data <= "110001000010";
      when "10101101100" => color_data <= "110101010010";
      when "10101101101" => color_data <= "101001000010";
      when "10101101110" => color_data <= "011000110010";
      when "10101101111" => color_data <= "110001000010";
      when "10101110000" => color_data <= "110001010010";
      when "10101110001" => color_data <= "110001000010";
      when "10101110010" => color_data <= "110001000010";
      when "10101110011" => color_data <= "110001000010";
      when "10101110100" => color_data <= "110001000010";
      when "10101110101" => color_data <= "110001000010";
      when "10101110110" => color_data <= "110001000010";
      when "10101110111" => color_data <= "110001000010";
      when "10101111000" => color_data <= "110001000010";
      when "10101111001" => color_data <= "110001000010";
      when "10101111010" => color_data <= "110001000010";
      when "10101111011" => color_data <= "110001000010";
      when "10101111100" => color_data <= "110001000010";
      when "10101111101" => color_data <= "110001000010";
      when "10101111110" => color_data <= "110001000010";
      when "10101111111" => color_data <= "110001010010";
      when "10110000000" => color_data <= "110101010010";
      when "10110000001" => color_data <= "110001010010";
      when "10110000010" => color_data <= "110001010010";
      when "10110000011" => color_data <= "110001010010";
      when "10110000100" => color_data <= "110001010010";
      when "10110000101" => color_data <= "110001010010";
      when "10110000110" => color_data <= "110001010010";
      when "10110000111" => color_data <= "111001010010";
      when "10110001000" => color_data <= "100001000010";
      when "10110001001" => color_data <= "011100110010";
      when "10110001010" => color_data <= "110101010010";
      when "10110001011" => color_data <= "110101010010";
      when "10110001100" => color_data <= "110001010010";
      when "10110001101" => color_data <= "110001010010";
      when "10110001110" => color_data <= "110001010010";
      when "10110001111" => color_data <= "110001010010";
      when "10110010000" => color_data <= "110001010010";
      when "10110010001" => color_data <= "110001010010";
      when "10110010010" => color_data <= "110001010010";
      when "10110010011" => color_data <= "110001010010";
      when "10110010100" => color_data <= "110001010010";
      when "10110010101" => color_data <= "110001010010";
      when "10110010110" => color_data <= "110001010010";
      when "10110010111" => color_data <= "110001010010";
      when "10110011000" => color_data <= "110001010010";
      when "10110011001" => color_data <= "110101010010";
      when "10110011010" => color_data <= "110101010010";
      when "10110011011" => color_data <= "011100110010";
      when "10110011100" => color_data <= "101001000010";
      when "10110011101" => color_data <= "111001010010";
      when "10110011110" => color_data <= "110001010010";
      when "10110011111" => color_data <= "110001010010";
      when "10110100000" => color_data <= "110001010010";
      when "10110100001" => color_data <= "110001010010";
      when "10110100010" => color_data <= "110001010010";
      when "10110100011" => color_data <= "110001010010";
      when "10110100100" => color_data <= "110001010010";
      when "10110100101" => color_data <= "110001010010";
      when "10110100110" => color_data <= "110001010010";
      when "10110100111" => color_data <= "110001010010";
      when "10110101000" => color_data <= "110001010010";
      when "10110101001" => color_data <= "110001010010";
      when "10110101010" => color_data <= "110001010010";
      when "10110101011" => color_data <= "110001010010";
      when "10110101100" => color_data <= "110101010010";
      when "10110101101" => color_data <= "101001000010";
      when "10110101110" => color_data <= "011000110010";
      when "10110101111" => color_data <= "110001010010";
      when "10110110000" => color_data <= "110101010010";
      when "10110110001" => color_data <= "110001010010";
      when "10110110010" => color_data <= "110001010010";
      when "10110110011" => color_data <= "110001010010";
      when "10110110100" => color_data <= "110001010010";
      when "10110110101" => color_data <= "110001010010";
      when "10110110110" => color_data <= "110001010010";
      when "10110110111" => color_data <= "110001010010";
      when "10110111000" => color_data <= "110001010010";
      when "10110111001" => color_data <= "110001010010";
      when "10110111010" => color_data <= "110001010010";
      when "10110111011" => color_data <= "110001010010";
      when "10110111100" => color_data <= "110001010010";
      when "10110111101" => color_data <= "110001010010";
      when "10110111110" => color_data <= "110001010010";
      when "10110111111" => color_data <= "110101010010";
      when "10111000000" => color_data <= "101001010010";
      when "10111000001" => color_data <= "101101000010";
      when "10111000010" => color_data <= "101001000010";
      when "10111000011" => color_data <= "101001000010";
      when "10111000100" => color_data <= "101001000010";
      when "10111000101" => color_data <= "101001000010";
      when "10111000110" => color_data <= "101001000010";
      when "10111000111" => color_data <= "101001000010";
      when "10111001000" => color_data <= "011100110010";
      when "10111001001" => color_data <= "011000110010";
      when "10111001010" => color_data <= "101001000010";
      when "10111001011" => color_data <= "101001000010";
      when "10111001100" => color_data <= "101001000010";
      when "10111001101" => color_data <= "101001000010";
      when "10111001110" => color_data <= "101001000010";
      when "10111001111" => color_data <= "101001000010";
      when "10111010000" => color_data <= "101001000010";
      when "10111010001" => color_data <= "101001000010";
      when "10111010010" => color_data <= "100101000010";
      when "10111010011" => color_data <= "101001000010";
      when "10111010100" => color_data <= "101001000010";
      when "10111010101" => color_data <= "100101000010";
      when "10111010110" => color_data <= "101001000010";
      when "10111010111" => color_data <= "101001000010";
      when "10111011000" => color_data <= "101001000010";
      when "10111011001" => color_data <= "101001000010";
      when "10111011010" => color_data <= "101001000010";
      when "10111011011" => color_data <= "010100110010";
      when "10111011100" => color_data <= "100000110010";
      when "10111011101" => color_data <= "101001000010";
      when "10111011110" => color_data <= "101001000010";
      when "10111011111" => color_data <= "101001000010";
      when "10111100000" => color_data <= "101001000010";
      when "10111100001" => color_data <= "101001000010";
      when "10111100010" => color_data <= "101001000010";
      when "10111100011" => color_data <= "101001000010";
      when "10111100100" => color_data <= "101001000010";
      when "10111100101" => color_data <= "101001000010";
      when "10111100110" => color_data <= "101001000010";
      when "10111100111" => color_data <= "101001000010";
      when "10111101000" => color_data <= "100101000010";
      when "10111101001" => color_data <= "101001000010";
      when "10111101010" => color_data <= "101001000010";
      when "10111101011" => color_data <= "101001000010";
      when "10111101100" => color_data <= "101001000010";
      when "10111101101" => color_data <= "100001000010";
      when "10111101110" => color_data <= "010100110010";
      when "10111101111" => color_data <= "101001000010";
      when "10111110000" => color_data <= "101001000010";
      when "10111110001" => color_data <= "101001000010";
      when "10111110010" => color_data <= "101001000010";
      when "10111110011" => color_data <= "101001000010";
      when "10111110100" => color_data <= "101001000010";
      when "10111110101" => color_data <= "101001000010";
      when "10111110110" => color_data <= "101001000010";
      when "10111110111" => color_data <= "100101000010";
      when "10111111000" => color_data <= "101001000010";
      when "10111111001" => color_data <= "101001000010";
      when "10111111010" => color_data <= "101001000010";
      when "10111111011" => color_data <= "101001000010";
      when "10111111100" => color_data <= "101001000010";
      when "10111111101" => color_data <= "101001000010";
      when "10111111110" => color_data <= "101001000010";
      when "10111111111" => color_data <= "101001010010";
      when "11000000000" => color_data <= "011101000010";
      when "11000000001" => color_data <= "010100110010";
      when "11000000010" => color_data <= "011100110010";
      when "11000000011" => color_data <= "011100110010";
      when "11000000100" => color_data <= "011100110010";
      when "11000000101" => color_data <= "011100110010";
      when "11000000110" => color_data <= "011100110010";
      when "11000000111" => color_data <= "011100110010";
      when "11000001000" => color_data <= "011100110010";
      when "11000001001" => color_data <= "100000110010";
      when "11000001010" => color_data <= "011100110010";
      when "11000001011" => color_data <= "011100110010";
      when "11000001100" => color_data <= "011100110010";
      when "11000001101" => color_data <= "011100110010";
      when "11000001110" => color_data <= "011100110010";
      when "11000001111" => color_data <= "011100110010";
      when "11000010000" => color_data <= "011100110010";
      when "11000010001" => color_data <= "011100110010";
      when "11000010010" => color_data <= "100000110010";
      when "11000010011" => color_data <= "011000110010";
      when "11000010100" => color_data <= "011000110010";
      when "11000010101" => color_data <= "100000110010";
      when "11000010110" => color_data <= "011100110010";
      when "11000010111" => color_data <= "011100110010";
      when "11000011000" => color_data <= "011100110010";
      when "11000011001" => color_data <= "011100110010";
      when "11000011010" => color_data <= "011100110010";
      when "11000011011" => color_data <= "100000110010";
      when "11000011100" => color_data <= "011100110010";
      when "11000011101" => color_data <= "011100110010";
      when "11000011110" => color_data <= "011100110010";
      when "11000011111" => color_data <= "011100110010";
      when "11000100000" => color_data <= "011100110010";
      when "11000100001" => color_data <= "011100110010";
      when "11000100010" => color_data <= "011100110010";
      when "11000100011" => color_data <= "011100110010";
      when "11000100100" => color_data <= "011100110010";
      when "11000100101" => color_data <= "011100110010";
      when "11000100110" => color_data <= "011000110010";
      when "11000100111" => color_data <= "011100110010";
      when "11000101000" => color_data <= "100000110010";
      when "11000101001" => color_data <= "011100110010";
      when "11000101010" => color_data <= "011100110010";
      when "11000101011" => color_data <= "011100110010";
      when "11000101100" => color_data <= "011100110010";
      when "11000101101" => color_data <= "011100110010";
      when "11000101110" => color_data <= "100000110010";
      when "11000101111" => color_data <= "011100110010";
      when "11000110000" => color_data <= "011100110010";
      when "11000110001" => color_data <= "011100110010";
      when "11000110010" => color_data <= "011100110010";
      when "11000110011" => color_data <= "011100110010";
      when "11000110100" => color_data <= "011100110010";
      when "11000110101" => color_data <= "011100110010";
      when "11000110110" => color_data <= "011100110010";
      when "11000110111" => color_data <= "100000110010";
      when "11000111000" => color_data <= "011100110010";
      when "11000111001" => color_data <= "011000110010";
      when "11000111010" => color_data <= "011100110010";
      when "11000111011" => color_data <= "011100110010";
      when "11000111100" => color_data <= "011100110010";
      when "11000111101" => color_data <= "011100110010";
      when "11000111110" => color_data <= "011100110010";
      when "11000111111" => color_data <= "100001000010";
      when "11001000000" => color_data <= "101101010010";
      when "11001000001" => color_data <= "011000110010";
      when "11001000010" => color_data <= "101101000010";
      when "11001000011" => color_data <= "110101010010";
      when "11001000100" => color_data <= "110001010010";
      when "11001000101" => color_data <= "110001010010";
      when "11001000110" => color_data <= "110001010010";
      when "11001000111" => color_data <= "110001010010";
      when "11001001000" => color_data <= "110001010010";
      when "11001001001" => color_data <= "110001010010";
      when "11001001010" => color_data <= "110001010010";
      when "11001001011" => color_data <= "110001010010";
      when "11001001100" => color_data <= "110001010010";
      when "11001001101" => color_data <= "110001010010";
      when "11001001110" => color_data <= "110001010010";
      when "11001001111" => color_data <= "110001010010";
      when "11001010000" => color_data <= "110001010010";
      when "11001010001" => color_data <= "110001010010";
      when "11001010010" => color_data <= "110101010010";
      when "11001010011" => color_data <= "100001000010";
      when "11001010100" => color_data <= "011100110010";
      when "11001010101" => color_data <= "110101010010";
      when "11001010110" => color_data <= "110001010010";
      when "11001010111" => color_data <= "110001010010";
      when "11001011000" => color_data <= "110001010010";
      when "11001011001" => color_data <= "110001010010";
      when "11001011010" => color_data <= "110001010010";
      when "11001011011" => color_data <= "110001010010";
      when "11001011100" => color_data <= "110001010010";
      when "11001011101" => color_data <= "110001010010";
      when "11001011110" => color_data <= "110001010010";
      when "11001011111" => color_data <= "110001010010";
      when "11001100000" => color_data <= "110001010010";
      when "11001100001" => color_data <= "110001010010";
      when "11001100010" => color_data <= "110001010010";
      when "11001100011" => color_data <= "110001010010";
      when "11001100100" => color_data <= "110001010010";
      when "11001100101" => color_data <= "110001010010";
      when "11001100110" => color_data <= "011000110010";
      when "11001100111" => color_data <= "101001000010";
      when "11001101000" => color_data <= "110101010010";
      when "11001101001" => color_data <= "110001010010";
      when "11001101010" => color_data <= "110001010010";
      when "11001101011" => color_data <= "110001010010";
      when "11001101100" => color_data <= "110001010010";
      when "11001101101" => color_data <= "110001010010";
      when "11001101110" => color_data <= "110001010010";
      when "11001101111" => color_data <= "110001010010";
      when "11001110000" => color_data <= "110001010010";
      when "11001110001" => color_data <= "110001010010";
      when "11001110010" => color_data <= "110001010010";
      when "11001110011" => color_data <= "110001010010";
      when "11001110100" => color_data <= "110001010010";
      when "11001110101" => color_data <= "110001010010";
      when "11001110110" => color_data <= "110001010010";
      when "11001110111" => color_data <= "110101010010";
      when "11001111000" => color_data <= "101001000010";
      when "11001111001" => color_data <= "011100110010";
      when "11001111010" => color_data <= "110101010010";
      when "11001111011" => color_data <= "110001010010";
      when "11001111100" => color_data <= "110001010010";
      when "11001111101" => color_data <= "110001010010";
      when "11001111110" => color_data <= "110001010010";
      when "11001111111" => color_data <= "110001010010";
      when "11010000000" => color_data <= "101101010010";
      when "11010000001" => color_data <= "011000110010";
      when "11010000010" => color_data <= "101101000010";
      when "11010000011" => color_data <= "110001010010";
      when "11010000100" => color_data <= "110001000010";
      when "11010000101" => color_data <= "110001000010";
      when "11010000110" => color_data <= "110001000010";
      when "11010000111" => color_data <= "110001000010";
      when "11010001000" => color_data <= "110001000010";
      when "11010001001" => color_data <= "110001000010";
      when "11010001010" => color_data <= "110001000010";
      when "11010001011" => color_data <= "110001000010";
      when "11010001100" => color_data <= "110001000010";
      when "11010001101" => color_data <= "110001000010";
      when "11010001110" => color_data <= "110001000010";
      when "11010001111" => color_data <= "110001000010";
      when "11010010000" => color_data <= "110001000010";
      when "11010010001" => color_data <= "110001000010";
      when "11010010010" => color_data <= "110101010010";
      when "11010010011" => color_data <= "100001000010";
      when "11010010100" => color_data <= "011100110010";
      when "11010010101" => color_data <= "110101010010";
      when "11010010110" => color_data <= "110001000010";
      when "11010010111" => color_data <= "110001000010";
      when "11010011000" => color_data <= "110001000010";
      when "11010011001" => color_data <= "110001000010";
      when "11010011010" => color_data <= "110001000010";
      when "11010011011" => color_data <= "110001000010";
      when "11010011100" => color_data <= "110001000010";
      when "11010011101" => color_data <= "110001000010";
      when "11010011110" => color_data <= "110001000010";
      when "11010011111" => color_data <= "110001000010";
      when "11010100000" => color_data <= "110001000010";
      when "11010100001" => color_data <= "110001000010";
      when "11010100010" => color_data <= "110001000010";
      when "11010100011" => color_data <= "110001000010";
      when "11010100100" => color_data <= "110001010010";
      when "11010100101" => color_data <= "110001010010";
      when "11010100110" => color_data <= "011000110010";
      when "11010100111" => color_data <= "101001000010";
      when "11010101000" => color_data <= "110101010010";
      when "11010101001" => color_data <= "110001000010";
      when "11010101010" => color_data <= "110001000010";
      when "11010101011" => color_data <= "110001000010";
      when "11010101100" => color_data <= "110001000010";
      when "11010101101" => color_data <= "110001000010";
      when "11010101110" => color_data <= "110001000010";
      when "11010101111" => color_data <= "110001000010";
      when "11010110000" => color_data <= "110001000010";
      when "11010110001" => color_data <= "110001000010";
      when "11010110010" => color_data <= "110001000010";
      when "11010110011" => color_data <= "110001000010";
      when "11010110100" => color_data <= "110001000010";
      when "11010110101" => color_data <= "110001000010";
      when "11010110110" => color_data <= "110001000010";
      when "11010110111" => color_data <= "110101010010";
      when "11010111000" => color_data <= "100101000010";
      when "11010111001" => color_data <= "011100110010";
      when "11010111010" => color_data <= "110001010010";
      when "11010111011" => color_data <= "110001000010";
      when "11010111100" => color_data <= "110001000010";
      when "11010111101" => color_data <= "110001000010";
      when "11010111110" => color_data <= "110001000010";
      when "11010111111" => color_data <= "110001010010";
      when "11011000000" => color_data <= "101101010010";
      when "11011000001" => color_data <= "011000110010";
      when "11011000010" => color_data <= "101101000010";
      when "11011000011" => color_data <= "110001010010";
      when "11011000100" => color_data <= "110001000010";
      when "11011000101" => color_data <= "110001000010";
      when "11011000110" => color_data <= "110001000010";
      when "11011000111" => color_data <= "110001000010";
      when "11011001000" => color_data <= "110001000010";
      when "11011001001" => color_data <= "110001000010";
      when "11011001010" => color_data <= "110001000010";
      when "11011001011" => color_data <= "110001000010";
      when "11011001100" => color_data <= "110001000010";
      when "11011001101" => color_data <= "110001000010";
      when "11011001110" => color_data <= "110001000010";
      when "11011001111" => color_data <= "110001000010";
      when "11011010000" => color_data <= "110001000010";
      when "11011010001" => color_data <= "110001000010";
      when "11011010010" => color_data <= "110101010010";
      when "11011010011" => color_data <= "100001000010";
      when "11011010100" => color_data <= "011100110010";
      when "11011010101" => color_data <= "110101010010";
      when "11011010110" => color_data <= "110001000010";
      when "11011010111" => color_data <= "110001000010";
      when "11011011000" => color_data <= "110001000010";
      when "11011011001" => color_data <= "110001000010";
      when "11011011010" => color_data <= "110001000010";
      when "11011011011" => color_data <= "110001000010";
      when "11011011100" => color_data <= "110001000010";
      when "11011011101" => color_data <= "110001000010";
      when "11011011110" => color_data <= "110001000010";
      when "11011011111" => color_data <= "110001000010";
      when "11011100000" => color_data <= "110001000010";
      when "11011100001" => color_data <= "110001000010";
      when "11011100010" => color_data <= "110001000010";
      when "11011100011" => color_data <= "110001000010";
      when "11011100100" => color_data <= "110001010010";
      when "11011100101" => color_data <= "110001010010";
      when "11011100110" => color_data <= "011000110010";
      when "11011100111" => color_data <= "100101000010";
      when "11011101000" => color_data <= "110101010010";
      when "11011101001" => color_data <= "110001000010";
      when "11011101010" => color_data <= "110001000010";
      when "11011101011" => color_data <= "110001000010";
      when "11011101100" => color_data <= "110001000010";
      when "11011101101" => color_data <= "110001000010";
      when "11011101110" => color_data <= "110001000010";
      when "11011101111" => color_data <= "110001000010";
      when "11011110000" => color_data <= "110001000010";
      when "11011110001" => color_data <= "110001000010";
      when "11011110010" => color_data <= "110001000010";
      when "11011110011" => color_data <= "110001000010";
      when "11011110100" => color_data <= "110001000010";
      when "11011110101" => color_data <= "110001000010";
      when "11011110110" => color_data <= "110001000010";
      when "11011110111" => color_data <= "110101010010";
      when "11011111000" => color_data <= "100101000010";
      when "11011111001" => color_data <= "011100110010";
      when "11011111010" => color_data <= "110001010010";
      when "11011111011" => color_data <= "110001000010";
      when "11011111100" => color_data <= "110001000010";
      when "11011111101" => color_data <= "110001000010";
      when "11011111110" => color_data <= "110001000010";
      when "11011111111" => color_data <= "110001010010";
      when "11100000000" => color_data <= "101101010010";
      when "11100000001" => color_data <= "011000110010";
      when "11100000010" => color_data <= "101101000010";
      when "11100000011" => color_data <= "110001010010";
      when "11100000100" => color_data <= "110001000010";
      when "11100000101" => color_data <= "110001000010";
      when "11100000110" => color_data <= "110001000010";
      when "11100000111" => color_data <= "110001000010";
      when "11100001000" => color_data <= "110001000010";
      when "11100001001" => color_data <= "110001000010";
      when "11100001010" => color_data <= "110001000010";
      when "11100001011" => color_data <= "110001000010";
      when "11100001100" => color_data <= "110001000010";
      when "11100001101" => color_data <= "110001000010";
      when "11100001110" => color_data <= "110001000010";
      when "11100001111" => color_data <= "110001000010";
      when "11100010000" => color_data <= "110001000010";
      when "11100010001" => color_data <= "110001000010";
      when "11100010010" => color_data <= "110101010010";
      when "11100010011" => color_data <= "100001000010";
      when "11100010100" => color_data <= "011100110010";
      when "11100010101" => color_data <= "110101010010";
      when "11100010110" => color_data <= "110001000010";
      when "11100010111" => color_data <= "110001000010";
      when "11100011000" => color_data <= "110001000010";
      when "11100011001" => color_data <= "110001000010";
      when "11100011010" => color_data <= "110001000010";
      when "11100011011" => color_data <= "110001000010";
      when "11100011100" => color_data <= "110001000010";
      when "11100011101" => color_data <= "110001000010";
      when "11100011110" => color_data <= "110001000010";
      when "11100011111" => color_data <= "110001000010";
      when "11100100000" => color_data <= "110001000010";
      when "11100100001" => color_data <= "110001000010";
      when "11100100010" => color_data <= "110001000010";
      when "11100100011" => color_data <= "110001000010";
      when "11100100100" => color_data <= "110001010010";
      when "11100100101" => color_data <= "110001010010";
      when "11100100110" => color_data <= "011000110010";
      when "11100100111" => color_data <= "100101000010";
      when "11100101000" => color_data <= "110101010010";
      when "11100101001" => color_data <= "110001000010";
      when "11100101010" => color_data <= "110001000010";
      when "11100101011" => color_data <= "110001000010";
      when "11100101100" => color_data <= "110001000010";
      when "11100101101" => color_data <= "110001000010";
      when "11100101110" => color_data <= "110001000010";
      when "11100101111" => color_data <= "110001000010";
      when "11100110000" => color_data <= "110001000010";
      when "11100110001" => color_data <= "110001000010";
      when "11100110010" => color_data <= "110001000010";
      when "11100110011" => color_data <= "110001000010";
      when "11100110100" => color_data <= "110001000010";
      when "11100110101" => color_data <= "110001000010";
      when "11100110110" => color_data <= "110001000010";
      when "11100110111" => color_data <= "110101010010";
      when "11100111000" => color_data <= "100101000010";
      when "11100111001" => color_data <= "011100110010";
      when "11100111010" => color_data <= "110001010010";
      when "11100111011" => color_data <= "110001000010";
      when "11100111100" => color_data <= "110001000010";
      when "11100111101" => color_data <= "110001000010";
      when "11100111110" => color_data <= "110001000010";
      when "11100111111" => color_data <= "110001010010";
      when "11101000000" => color_data <= "101101010010";
      when "11101000001" => color_data <= "011000110010";
      when "11101000010" => color_data <= "101101000010";
      when "11101000011" => color_data <= "110001010010";
      when "11101000100" => color_data <= "110001000010";
      when "11101000101" => color_data <= "110001000010";
      when "11101000110" => color_data <= "110001000010";
      when "11101000111" => color_data <= "110001000010";
      when "11101001000" => color_data <= "110001000010";
      when "11101001001" => color_data <= "110001000010";
      when "11101001010" => color_data <= "110001000010";
      when "11101001011" => color_data <= "110001000010";
      when "11101001100" => color_data <= "110001000010";
      when "11101001101" => color_data <= "110001000010";
      when "11101001110" => color_data <= "110001000010";
      when "11101001111" => color_data <= "110001000010";
      when "11101010000" => color_data <= "110001000010";
      when "11101010001" => color_data <= "110001000010";
      when "11101010010" => color_data <= "110101010010";
      when "11101010011" => color_data <= "100001000010";
      when "11101010100" => color_data <= "011100110010";
      when "11101010101" => color_data <= "110101010010";
      when "11101010110" => color_data <= "110001000010";
      when "11101010111" => color_data <= "110001000010";
      when "11101011000" => color_data <= "110001000010";
      when "11101011001" => color_data <= "110001000010";
      when "11101011010" => color_data <= "110001000010";
      when "11101011011" => color_data <= "110001000010";
      when "11101011100" => color_data <= "110001000010";
      when "11101011101" => color_data <= "110001000010";
      when "11101011110" => color_data <= "110001000010";
      when "11101011111" => color_data <= "110001000010";
      when "11101100000" => color_data <= "110001000010";
      when "11101100001" => color_data <= "110001000010";
      when "11101100010" => color_data <= "110001000010";
      when "11101100011" => color_data <= "110001000010";
      when "11101100100" => color_data <= "110001010010";
      when "11101100101" => color_data <= "110001010010";
      when "11101100110" => color_data <= "011000110010";
      when "11101100111" => color_data <= "100101000010";
      when "11101101000" => color_data <= "110101010010";
      when "11101101001" => color_data <= "110001000010";
      when "11101101010" => color_data <= "110001000010";
      when "11101101011" => color_data <= "110001000010";
      when "11101101100" => color_data <= "110001000010";
      when "11101101101" => color_data <= "110001000010";
      when "11101101110" => color_data <= "110001000010";
      when "11101101111" => color_data <= "110001000010";
      when "11101110000" => color_data <= "110001000010";
      when "11101110001" => color_data <= "110001000010";
      when "11101110010" => color_data <= "110001000010";
      when "11101110011" => color_data <= "110001000010";
      when "11101110100" => color_data <= "110001000010";
      when "11101110101" => color_data <= "110001000010";
      when "11101110110" => color_data <= "110001000010";
      when "11101110111" => color_data <= "110101010010";
      when "11101111000" => color_data <= "100101000010";
      when "11101111001" => color_data <= "011100110010";
      when "11101111010" => color_data <= "110001010010";
      when "11101111011" => color_data <= "110001000010";
      when "11101111100" => color_data <= "110001000010";
      when "11101111101" => color_data <= "110001000010";
      when "11101111110" => color_data <= "110001000010";
      when "11101111111" => color_data <= "110001010010";
      when "11110000000" => color_data <= "101101010010";
      when "11110000001" => color_data <= "011000110010";
      when "11110000010" => color_data <= "101101000010";
      when "11110000011" => color_data <= "110001010010";
      when "11110000100" => color_data <= "110001000010";
      when "11110000101" => color_data <= "110001000010";
      when "11110000110" => color_data <= "110001000010";
      when "11110000111" => color_data <= "110001000010";
      when "11110001000" => color_data <= "110001000010";
      when "11110001001" => color_data <= "110001000010";
      when "11110001010" => color_data <= "110001000010";
      when "11110001011" => color_data <= "110001000010";
      when "11110001100" => color_data <= "110001000010";
      when "11110001101" => color_data <= "110001000010";
      when "11110001110" => color_data <= "110001000010";
      when "11110001111" => color_data <= "110001000010";
      when "11110010000" => color_data <= "110001000010";
      when "11110010001" => color_data <= "110001000010";
      when "11110010010" => color_data <= "110101010010";
      when "11110010011" => color_data <= "100001000010";
      when "11110010100" => color_data <= "011100110010";
      when "11110010101" => color_data <= "110101010010";
      when "11110010110" => color_data <= "110001000010";
      when "11110010111" => color_data <= "110001000010";
      when "11110011000" => color_data <= "110001000010";
      when "11110011001" => color_data <= "110001000010";
      when "11110011010" => color_data <= "110001000010";
      when "11110011011" => color_data <= "110001000010";
      when "11110011100" => color_data <= "110001000010";
      when "11110011101" => color_data <= "110001000010";
      when "11110011110" => color_data <= "110001000010";
      when "11110011111" => color_data <= "110001000010";
      when "11110100000" => color_data <= "110001000010";
      when "11110100001" => color_data <= "110001000010";
      when "11110100010" => color_data <= "110001000010";
      when "11110100011" => color_data <= "110001000010";
      when "11110100100" => color_data <= "110001010010";
      when "11110100101" => color_data <= "110001010010";
      when "11110100110" => color_data <= "011000110010";
      when "11110100111" => color_data <= "100101000010";
      when "11110101000" => color_data <= "110101010010";
      when "11110101001" => color_data <= "110001000010";
      when "11110101010" => color_data <= "110001000010";
      when "11110101011" => color_data <= "110001000010";
      when "11110101100" => color_data <= "110001000010";
      when "11110101101" => color_data <= "110001000010";
      when "11110101110" => color_data <= "110001000010";
      when "11110101111" => color_data <= "110001000010";
      when "11110110000" => color_data <= "110001000010";
      when "11110110001" => color_data <= "110001000010";
      when "11110110010" => color_data <= "110001000010";
      when "11110110011" => color_data <= "110001000010";
      when "11110110100" => color_data <= "110001000010";
      when "11110110101" => color_data <= "110001000010";
      when "11110110110" => color_data <= "110001000010";
      when "11110110111" => color_data <= "110101010010";
      when "11110111000" => color_data <= "100101000010";
      when "11110111001" => color_data <= "011100110010";
      when "11110111010" => color_data <= "110001010010";
      when "11110111011" => color_data <= "110001000010";
      when "11110111100" => color_data <= "110001000010";
      when "11110111101" => color_data <= "110001000010";
      when "11110111110" => color_data <= "110001000010";
      when "11110111111" => color_data <= "110001010010";
      when "11111000000" => color_data <= "101101010011";
      when "11111000001" => color_data <= "011000110010";
      when "11111000010" => color_data <= "101101010010";
      when "11111000011" => color_data <= "110001010010";
      when "11111000100" => color_data <= "110001010010";
      when "11111000101" => color_data <= "110001010010";
      when "11111000110" => color_data <= "110001010010";
      when "11111000111" => color_data <= "110001010010";
      when "11111001000" => color_data <= "110001010010";
      when "11111001001" => color_data <= "110001010010";
      when "11111001010" => color_data <= "110001010010";
      when "11111001011" => color_data <= "110001010010";
      when "11111001100" => color_data <= "110001010010";
      when "11111001101" => color_data <= "110001010010";
      when "11111001110" => color_data <= "110001010010";
      when "11111001111" => color_data <= "110001010010";
      when "11111010000" => color_data <= "110001010010";
      when "11111010001" => color_data <= "110001010010";
      when "11111010010" => color_data <= "110101010010";
      when "11111010011" => color_data <= "100101000010";
      when "11111010100" => color_data <= "011101000010";
      when "11111010101" => color_data <= "110101010010";
      when "11111010110" => color_data <= "110001010010";
      when "11111010111" => color_data <= "110001010010";
      when "11111011000" => color_data <= "110001010010";
      when "11111011001" => color_data <= "110001010010";
      when "11111011010" => color_data <= "110001010010";
      when "11111011011" => color_data <= "110001010010";
      when "11111011100" => color_data <= "110001010010";
      when "11111011101" => color_data <= "110001010010";
      when "11111011110" => color_data <= "110001010010";
      when "11111011111" => color_data <= "110001010010";
      when "11111100000" => color_data <= "110001010010";
      when "11111100001" => color_data <= "110001010010";
      when "11111100010" => color_data <= "110001010010";
      when "11111100011" => color_data <= "110001010010";
      when "11111100100" => color_data <= "110001010010";
      when "11111100101" => color_data <= "110001010010";
      when "11111100110" => color_data <= "011101000010";
      when "11111100111" => color_data <= "101001000010";
      when "11111101000" => color_data <= "110101010010";
      when "11111101001" => color_data <= "110001010010";
      when "11111101010" => color_data <= "110001010010";
      when "11111101011" => color_data <= "110001010010";
      when "11111101100" => color_data <= "110001010010";
      when "11111101101" => color_data <= "110001010010";
      when "11111101110" => color_data <= "110001010010";
      when "11111101111" => color_data <= "110001010010";
      when "11111110000" => color_data <= "110001010010";
      when "11111110001" => color_data <= "110001010010";
      when "11111110010" => color_data <= "110001010010";
      when "11111110011" => color_data <= "110001010010";
      when "11111110100" => color_data <= "110001010010";
      when "11111110101" => color_data <= "110001010010";
      when "11111110110" => color_data <= "110001010010";
      when "11111110111" => color_data <= "110101010010";
      when "11111111000" => color_data <= "101001000010";
      when "11111111001" => color_data <= "011101000010";
      when "11111111010" => color_data <= "110001010010";
      when "11111111011" => color_data <= "110001010010";
      when "11111111100" => color_data <= "110001010010";
      when "11111111101" => color_data <= "110001010010";
      when "11111111110" => color_data <= "110001000010";
      when "11111111111" => color_data <= "110001100011";
      when others => color_data <= (others => '0');
    end case;
  end process;
end Behavioral;
