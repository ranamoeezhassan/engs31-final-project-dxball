library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity paddle_rom is
  Port (
    clk        : in  std_logic;
    row        : in  std_logic_vector(3 downto 0);
    col        : in  std_logic_vector(6 downto 0);
    color_data : out std_logic_vector(11 downto 0)
  );
end entity;

architecture Behavioral of paddle_rom is
  signal addr : std_logic_vector(10 downto 0);
  signal row_reg : std_logic_vector(3 downto 0);
  signal col_reg : std_logic_vector(6 downto 0);
begin

  process(clk)
  begin
    if rising_edge(clk) then
      row_reg <= row;
      col_reg <= col;
    end if;
  end process;

  addr <= row_reg & col_reg;

  process(addr)
  begin
    case addr is
      when "00000000000" => color_data <= "000000000000";
      when "00000000001" => color_data <= "000000000000";
      when "00000000010" => color_data <= "000000000000";
      when "00000000011" => color_data <= "000000000000";
      when "00000000100" => color_data <= "000000000000";
      when "00000000101" => color_data <= "000000000000";
      when "00000000110" => color_data <= "000000000000";
      when "00000000111" => color_data <= "000000000000";
      when "00000001000" => color_data <= "000000000000";
      when "00000001001" => color_data <= "000000000000";
      when "00000001010" => color_data <= "000000000000";
      when "00000001011" => color_data <= "000000000000";
      when "00000001100" => color_data <= "000000000000";
      when "00000001101" => color_data <= "000000000000";
      when "00000001110" => color_data <= "000000000000";
      when "00000001111" => color_data <= "000000000000";
      when "00000010000" => color_data <= "000000000000";
      when "00000010001" => color_data <= "000000000000";
      when "00000010010" => color_data <= "000000000000";
      when "00000010011" => color_data <= "000000000000";
      when "00000010100" => color_data <= "000000000000";
      when "00000010101" => color_data <= "000000000000";
      when "00000010110" => color_data <= "000000000000";
      when "00000010111" => color_data <= "000000000000";
      when "00000011000" => color_data <= "000000000000";
      when "00000011001" => color_data <= "000000000000";
      when "00000011010" => color_data <= "000000000000";
      when "00000011011" => color_data <= "000000000000";
      when "00000011100" => color_data <= "000000000000";
      when "00000011101" => color_data <= "000000000000";
      when "00000011110" => color_data <= "000000000000";
      when "00000011111" => color_data <= "000000000000";
      when "00000100000" => color_data <= "000000000000";
      when "00000100001" => color_data <= "000000000000";
      when "00000100010" => color_data <= "000000000000";
      when "00000100011" => color_data <= "000000000000";
      when "00000100100" => color_data <= "000000000000";
      when "00000100101" => color_data <= "000000000000";
      when "00000100110" => color_data <= "000000000000";
      when "00000100111" => color_data <= "000000000000";
      when "00000101000" => color_data <= "000000000000";
      when "00000101001" => color_data <= "000000000000";
      when "00000101010" => color_data <= "000000000000";
      when "00000101011" => color_data <= "000000000000";
      when "00000101100" => color_data <= "000000000000";
      when "00000101101" => color_data <= "000000000000";
      when "00000101110" => color_data <= "000100010000";
      when "00000101111" => color_data <= "000100010000";
      when "00000110000" => color_data <= "000100010000";
      when "00000110001" => color_data <= "001000010000";
      when "00000110010" => color_data <= "001100100001";
      when "00000110011" => color_data <= "001100110001";
      when "00000110100" => color_data <= "010000110001";
      when "00000110101" => color_data <= "010000110001";
      when "00000110110" => color_data <= "010101000001";
      when "00000110111" => color_data <= "010101000010";
      when "00000111000" => color_data <= "010101000001";
      when "00000111001" => color_data <= "011001010010";
      when "00000111010" => color_data <= "011101100011";
      when "00000111011" => color_data <= "011101010010";
      when "00000111100" => color_data <= "011101100010";
      when "00000111101" => color_data <= "100001100010";
      when "00000111110" => color_data <= "100001100011";
      when "00000111111" => color_data <= "100101110011";
      when "00001000000" => color_data <= "100101110010";
      when "00001000001" => color_data <= "100101110010";
      when "00001000010" => color_data <= "101010000011";
      when "00001000011" => color_data <= "101110000011";
      when "00001000100" => color_data <= "101110000011";
      when "00001000101" => color_data <= "110010010100";
      when "00001000110" => color_data <= "110110100100";
      when "00001000111" => color_data <= "110110100100";
      when "00001001000" => color_data <= "111010110100";
      when "00001001001" => color_data <= "111111000101";
      when "00001001010" => color_data <= "111111000100";
      when "00001001011" => color_data <= "111111000100";
      when "00001001100" => color_data <= "111010110100";
      when "00001001101" => color_data <= "100110000011";
      when "00001001110" => color_data <= "000100000000";
      when "00001001111" => color_data <= "000000000000";
      when "00010000000" => color_data <= "000000000000";
      when "00010000001" => color_data <= "000000000000";
      when "00010000010" => color_data <= "000000000000";
      when "00010000011" => color_data <= "000000000000";
      when "00010000100" => color_data <= "000000000000";
      when "00010000101" => color_data <= "000000000000";
      when "00010000110" => color_data <= "000000000000";
      when "00010000111" => color_data <= "000000000000";
      when "00010001000" => color_data <= "000000000000";
      when "00010001001" => color_data <= "000000000000";
      when "00010001010" => color_data <= "000000000000";
      when "00010001011" => color_data <= "000000000000";
      when "00010001100" => color_data <= "000000000000";
      when "00010001101" => color_data <= "000000000000";
      when "00010001110" => color_data <= "000000000000";
      when "00010001111" => color_data <= "000000000000";
      when "00010010000" => color_data <= "000000000000";
      when "00010010001" => color_data <= "000000000000";
      when "00010010010" => color_data <= "000000000000";
      when "00010010011" => color_data <= "000000000000";
      when "00010010100" => color_data <= "000000000000";
      when "00010010101" => color_data <= "000000000000";
      when "00010010110" => color_data <= "000000000000";
      when "00010010111" => color_data <= "000000000000";
      when "00010011000" => color_data <= "000000000000";
      when "00010011001" => color_data <= "000000000000";
      when "00010011010" => color_data <= "000000000000";
      when "00010011011" => color_data <= "000000000000";
      when "00010011100" => color_data <= "000000000000";
      when "00010011101" => color_data <= "000000000000";
      when "00010011110" => color_data <= "000000000000";
      when "00010011111" => color_data <= "000000000000";
      when "00010100000" => color_data <= "000000000000";
      when "00010100001" => color_data <= "000000000000";
      when "00010100010" => color_data <= "000000000000";
      when "00010100011" => color_data <= "000000000000";
      when "00010100100" => color_data <= "000000000000";
      when "00010100101" => color_data <= "000000000000";
      when "00010100110" => color_data <= "000000000000";
      when "00010100111" => color_data <= "001000100001";
      when "00010101000" => color_data <= "010101000001";
      when "00010101001" => color_data <= "011101100010";
      when "00010101010" => color_data <= "101010000011";
      when "00010101011" => color_data <= "110010010011";
      when "00010101100" => color_data <= "110110100100";
      when "00010101101" => color_data <= "111010110100";
      when "00010101110" => color_data <= "111110110100";
      when "00010101111" => color_data <= "111111000100";
      when "00010110000" => color_data <= "111111000100";
      when "00010110001" => color_data <= "111111000100";
      when "00010110010" => color_data <= "111111010101";
      when "00010110011" => color_data <= "111111010101";
      when "00010110100" => color_data <= "111111010100";
      when "00010110101" => color_data <= "111111010100";
      when "00010110110" => color_data <= "111111010101";
      when "00010110111" => color_data <= "111111010101";
      when "00010111000" => color_data <= "111111010101";
      when "00010111001" => color_data <= "111111100101";
      when "00010111010" => color_data <= "111111100101";
      when "00010111011" => color_data <= "111111100101";
      when "00010111100" => color_data <= "111111100101";
      when "00010111101" => color_data <= "111111100101";
      when "00010111110" => color_data <= "111111100101";
      when "00010111111" => color_data <= "111111100101";
      when "00011000000" => color_data <= "111111100101";
      when "00011000001" => color_data <= "111111100101";
      when "00011000010" => color_data <= "111111010101";
      when "00011000011" => color_data <= "111111010101";
      when "00011000100" => color_data <= "111111010101";
      when "00011000101" => color_data <= "111111010100";
      when "00011000110" => color_data <= "111111000100";
      when "00011000111" => color_data <= "111111000100";
      when "00011001000" => color_data <= "111111000100";
      when "00011001001" => color_data <= "111110110011";
      when "00011001010" => color_data <= "111110110100";
      when "00011001011" => color_data <= "111110110100";
      when "00011001100" => color_data <= "111111000100";
      when "00011001101" => color_data <= "111111110101";
      when "00011001110" => color_data <= "111010110100";
      when "00011001111" => color_data <= "000000000000";
      when "00100000000" => color_data <= "000000000000";
      when "00100000001" => color_data <= "000100010001";
      when "00100000010" => color_data <= "000100010000";
      when "00100000011" => color_data <= "000000000000";
      when "00100000100" => color_data <= "000000000000";
      when "00100000101" => color_data <= "000000000000";
      when "00100000110" => color_data <= "000000000000";
      when "00100000111" => color_data <= "000000000000";
      when "00100001000" => color_data <= "000000000000";
      when "00100001001" => color_data <= "000000000000";
      when "00100001010" => color_data <= "000000000000";
      when "00100001011" => color_data <= "000000000000";
      when "00100001100" => color_data <= "000000000000";
      when "00100001101" => color_data <= "000000000000";
      when "00100001110" => color_data <= "000000000000";
      when "00100001111" => color_data <= "000000000000";
      when "00100010000" => color_data <= "000000000000";
      when "00100010001" => color_data <= "000000000000";
      when "00100010010" => color_data <= "000000000000";
      when "00100010011" => color_data <= "000000000000";
      when "00100010100" => color_data <= "000000000000";
      when "00100010101" => color_data <= "000000000000";
      when "00100010110" => color_data <= "000000000000";
      when "00100010111" => color_data <= "000000000000";
      when "00100011000" => color_data <= "000000000000";
      when "00100011001" => color_data <= "000000000000";
      when "00100011010" => color_data <= "000000000000";
      when "00100011011" => color_data <= "000000000000";
      when "00100011100" => color_data <= "000000000000";
      when "00100011101" => color_data <= "000000000000";
      when "00100011110" => color_data <= "000000000000";
      when "00100011111" => color_data <= "000000000000";
      when "00100100000" => color_data <= "000100010000";
      when "00100100001" => color_data <= "001100100001";
      when "00100100010" => color_data <= "011001010010";
      when "00100100011" => color_data <= "100101110011";
      when "00100100100" => color_data <= "101010000011";
      when "00100100101" => color_data <= "110010100100";
      when "00100100110" => color_data <= "111010110100";
      when "00100100111" => color_data <= "111111000100";
      when "00100101000" => color_data <= "111111010101";
      when "00100101001" => color_data <= "111111100101";
      when "00100101010" => color_data <= "111111100101";
      when "00100101011" => color_data <= "111111010100";
      when "00100101100" => color_data <= "111111010100";
      when "00100101101" => color_data <= "111111000100";
      when "00100101110" => color_data <= "111111000100";
      when "00100101111" => color_data <= "111111000100";
      when "00100110000" => color_data <= "111111000100";
      when "00100110001" => color_data <= "111111000100";
      when "00100110010" => color_data <= "111111000100";
      when "00100110011" => color_data <= "111111000100";
      when "00100110100" => color_data <= "111111000100";
      when "00100110101" => color_data <= "111111000100";
      when "00100110110" => color_data <= "111111000100";
      when "00100110111" => color_data <= "111111000100";
      when "00100111000" => color_data <= "111111000100";
      when "00100111001" => color_data <= "111111000100";
      when "00100111010" => color_data <= "111110110100";
      when "00100111011" => color_data <= "111110110100";
      when "00100111100" => color_data <= "111110110100";
      when "00100111101" => color_data <= "111110110100";
      when "00100111110" => color_data <= "111110110100";
      when "00100111111" => color_data <= "111110110100";
      when "00101000000" => color_data <= "111110110100";
      when "00101000001" => color_data <= "111110110100";
      when "00101000010" => color_data <= "111110110100";
      when "00101000011" => color_data <= "111110110100";
      when "00101000100" => color_data <= "111110110100";
      when "00101000101" => color_data <= "111110110100";
      when "00101000110" => color_data <= "111110110100";
      when "00101000111" => color_data <= "111110110100";
      when "00101001000" => color_data <= "111110110100";
      when "00101001001" => color_data <= "111110110100";
      when "00101001010" => color_data <= "111110110100";
      when "00101001011" => color_data <= "111110110100";
      when "00101001100" => color_data <= "111110110100";
      when "00101001101" => color_data <= "111110110100";
      when "00101001110" => color_data <= "111111110101";
      when "00101001111" => color_data <= "100001100010";
      when "00110000000" => color_data <= "010000110010";
      when "00110000001" => color_data <= "111111100111";
      when "00110000010" => color_data <= "111111010110";
      when "00110000011" => color_data <= "010101000010";
      when "00110000100" => color_data <= "001100110001";
      when "00110000101" => color_data <= "001000010001";
      when "00110000110" => color_data <= "000000000000";
      when "00110000111" => color_data <= "000000000000";
      when "00110001000" => color_data <= "000000000000";
      when "00110001001" => color_data <= "000000000000";
      when "00110001010" => color_data <= "000000000000";
      when "00110001011" => color_data <= "000000000000";
      when "00110001100" => color_data <= "000000000000";
      when "00110001101" => color_data <= "000000000000";
      when "00110001110" => color_data <= "000000000000";
      when "00110001111" => color_data <= "000000000000";
      when "00110010000" => color_data <= "000000000000";
      when "00110010001" => color_data <= "000000000000";
      when "00110010010" => color_data <= "000000000000";
      when "00110010011" => color_data <= "000000000000";
      when "00110010100" => color_data <= "000000000000";
      when "00110010101" => color_data <= "000000000000";
      when "00110010110" => color_data <= "000000000000";
      when "00110010111" => color_data <= "000000000000";
      when "00110011000" => color_data <= "000000000000";
      when "00110011001" => color_data <= "000000000000";
      when "00110011010" => color_data <= "000100010000";
      when "00110011011" => color_data <= "010101000010";
      when "00110011100" => color_data <= "011101100010";
      when "00110011101" => color_data <= "100101110011";
      when "00110011110" => color_data <= "101110010011";
      when "00110011111" => color_data <= "110110100100";
      when "00110100000" => color_data <= "111111000100";
      when "00110100001" => color_data <= "111111000100";
      when "00110100010" => color_data <= "111111010101";
      when "00110100011" => color_data <= "111111100101";
      when "00110100100" => color_data <= "111111010101";
      when "00110100101" => color_data <= "111111010100";
      when "00110100110" => color_data <= "111111000100";
      when "00110100111" => color_data <= "111111000100";
      when "00110101000" => color_data <= "111111000100";
      when "00110101001" => color_data <= "111110110100";
      when "00110101010" => color_data <= "111110110100";
      when "00110101011" => color_data <= "111110110100";
      when "00110101100" => color_data <= "111110110100";
      when "00110101101" => color_data <= "111110110100";
      when "00110101110" => color_data <= "111110110100";
      when "00110101111" => color_data <= "111110110100";
      when "00110110000" => color_data <= "111110110100";
      when "00110110001" => color_data <= "111110110100";
      when "00110110010" => color_data <= "111110110100";
      when "00110110011" => color_data <= "111110110100";
      when "00110110100" => color_data <= "111110110100";
      when "00110110101" => color_data <= "111110110100";
      when "00110110110" => color_data <= "111110110100";
      when "00110110111" => color_data <= "111110110100";
      when "00110111000" => color_data <= "111110110100";
      when "00110111001" => color_data <= "111110110100";
      when "00110111010" => color_data <= "111110110100";
      when "00110111011" => color_data <= "111110110100";
      when "00110111100" => color_data <= "111110110100";
      when "00110111101" => color_data <= "111110110100";
      when "00110111110" => color_data <= "111110110100";
      when "00110111111" => color_data <= "111110110100";
      when "00111000000" => color_data <= "111110110100";
      when "00111000001" => color_data <= "111110110100";
      when "00111000010" => color_data <= "111110110100";
      when "00111000011" => color_data <= "111110110100";
      when "00111000100" => color_data <= "111110110100";
      when "00111000101" => color_data <= "111110110100";
      when "00111000110" => color_data <= "111110110100";
      when "00111000111" => color_data <= "111110110100";
      when "00111001000" => color_data <= "111110110100";
      when "00111001001" => color_data <= "111110110100";
      when "00111001010" => color_data <= "111110110100";
      when "00111001011" => color_data <= "111110110100";
      when "00111001100" => color_data <= "111110110100";
      when "00111001101" => color_data <= "111110110100";
      when "00111001110" => color_data <= "111111010100";
      when "00111001111" => color_data <= "110010100011";
      when "01000000000" => color_data <= "110110110110";
      when "01000000001" => color_data <= "111111110111";
      when "01000000010" => color_data <= "111111010111";
      when "01000000011" => color_data <= "111111100110";
      when "01000000100" => color_data <= "111111100101";
      when "01000000101" => color_data <= "011101100011";
      when "01000000110" => color_data <= "000000010010";
      when "01000000111" => color_data <= "001000110011";
      when "01000001000" => color_data <= "001000110011";
      when "01000001001" => color_data <= "001000110011";
      when "01000001010" => color_data <= "001000110011";
      when "01000001011" => color_data <= "001000110011";
      when "01000001100" => color_data <= "001000110011";
      when "01000001101" => color_data <= "001000110011";
      when "01000001110" => color_data <= "001000110011";
      when "01000001111" => color_data <= "001000110011";
      when "01000010000" => color_data <= "001000110011";
      when "01000010001" => color_data <= "001000110011";
      when "01000010010" => color_data <= "001000110011";
      when "01000010011" => color_data <= "001000110011";
      when "01000010100" => color_data <= "001000110011";
      when "01000010101" => color_data <= "001000110011";
      when "01000010110" => color_data <= "001000110011";
      when "01000010111" => color_data <= "001000110011";
      when "01000011000" => color_data <= "001000110011";
      when "01000011001" => color_data <= "000000010011";
      when "01000011010" => color_data <= "011001010011";
      when "01000011011" => color_data <= "111111100101";
      when "01000011100" => color_data <= "111111100101";
      when "01000011101" => color_data <= "111111100101";
      when "01000011110" => color_data <= "111111010101";
      when "01000011111" => color_data <= "111111010100";
      when "01000100000" => color_data <= "111111000100";
      when "01000100001" => color_data <= "111111000100";
      when "01000100010" => color_data <= "111111000100";
      when "01000100011" => color_data <= "111110110100";
      when "01000100100" => color_data <= "111110110100";
      when "01000100101" => color_data <= "111110110100";
      when "01000100110" => color_data <= "111110110100";
      when "01000100111" => color_data <= "111110110100";
      when "01000101000" => color_data <= "111110110100";
      when "01000101001" => color_data <= "111110110100";
      when "01000101010" => color_data <= "111110110100";
      when "01000101011" => color_data <= "111110110100";
      when "01000101100" => color_data <= "111110110100";
      when "01000101101" => color_data <= "111110110100";
      when "01000101110" => color_data <= "111110110100";
      when "01000101111" => color_data <= "111110110100";
      when "01000110000" => color_data <= "111110110100";
      when "01000110001" => color_data <= "111110110100";
      when "01000110010" => color_data <= "111110110100";
      when "01000110011" => color_data <= "111110110100";
      when "01000110100" => color_data <= "111110110100";
      when "01000110101" => color_data <= "111110110100";
      when "01000110110" => color_data <= "111110110100";
      when "01000110111" => color_data <= "111110110100";
      when "01000111000" => color_data <= "111110110100";
      when "01000111001" => color_data <= "111110110100";
      when "01000111010" => color_data <= "111110110100";
      when "01000111011" => color_data <= "111110110100";
      when "01000111100" => color_data <= "111110110100";
      when "01000111101" => color_data <= "111110110100";
      when "01000111110" => color_data <= "111110110100";
      when "01000111111" => color_data <= "111110110100";
      when "01001000000" => color_data <= "111110110100";
      when "01001000001" => color_data <= "111110110100";
      when "01001000010" => color_data <= "111110110100";
      when "01001000011" => color_data <= "111110110100";
      when "01001000100" => color_data <= "111110110100";
      when "01001000101" => color_data <= "111110110100";
      when "01001000110" => color_data <= "111110110100";
      when "01001000111" => color_data <= "111110110100";
      when "01001001000" => color_data <= "111110110100";
      when "01001001001" => color_data <= "111110110100";
      when "01001001010" => color_data <= "111110110100";
      when "01001001011" => color_data <= "111110110100";
      when "01001001100" => color_data <= "111110110100";
      when "01001001101" => color_data <= "111110110100";
      when "01001001110" => color_data <= "111111010100";
      when "01001001111" => color_data <= "110110100100";
      when "01010000000" => color_data <= "111111000110";
      when "01010000001" => color_data <= "111111010110";
      when "01010000010" => color_data <= "111111010111";
      when "01010000011" => color_data <= "111111010110";
      when "01010000100" => color_data <= "111111000100";
      when "01010000101" => color_data <= "011001010011";
      when "01010000110" => color_data <= "000000010010";
      when "01010000111" => color_data <= "001000110011";
      when "01010001000" => color_data <= "001000110011";
      when "01010001001" => color_data <= "001000100011";
      when "01010001010" => color_data <= "001000110011";
      when "01010001011" => color_data <= "001000110011";
      when "01010001100" => color_data <= "001000100011";
      when "01010001101" => color_data <= "001000110011";
      when "01010001110" => color_data <= "001000110011";
      when "01010001111" => color_data <= "001000100011";
      when "01010010000" => color_data <= "001000100011";
      when "01010010001" => color_data <= "001000110011";
      when "01010010010" => color_data <= "001000100011";
      when "01010010011" => color_data <= "001000100011";
      when "01010010100" => color_data <= "001000110011";
      when "01010010101" => color_data <= "001000110011";
      when "01010010110" => color_data <= "001000100011";
      when "01010010111" => color_data <= "001000100011";
      when "01010011000" => color_data <= "001000100011";
      when "01010011001" => color_data <= "000000010010";
      when "01010011010" => color_data <= "010101010011";
      when "01010011011" => color_data <= "111111000100";
      when "01010011100" => color_data <= "111110110011";
      when "01010011101" => color_data <= "111110110100";
      when "01010011110" => color_data <= "111110110100";
      when "01010011111" => color_data <= "111110110100";
      when "01010100000" => color_data <= "111110110100";
      when "01010100001" => color_data <= "111110110100";
      when "01010100010" => color_data <= "111110110100";
      when "01010100011" => color_data <= "111111000100";
      when "01010100100" => color_data <= "111111000100";
      when "01010100101" => color_data <= "111111000100";
      when "01010100110" => color_data <= "111111000100";
      when "01010100111" => color_data <= "111111000100";
      when "01010101000" => color_data <= "111111000100";
      when "01010101001" => color_data <= "111111000100";
      when "01010101010" => color_data <= "111111000100";
      when "01010101011" => color_data <= "111111000100";
      when "01010101100" => color_data <= "111110110100";
      when "01010101101" => color_data <= "111110110100";
      when "01010101110" => color_data <= "111110110100";
      when "01010101111" => color_data <= "111110110100";
      when "01010110000" => color_data <= "111110110100";
      when "01010110001" => color_data <= "111110110100";
      when "01010110010" => color_data <= "111110110100";
      when "01010110011" => color_data <= "111110110100";
      when "01010110100" => color_data <= "111110110100";
      when "01010110101" => color_data <= "111110110100";
      when "01010110110" => color_data <= "111110110100";
      when "01010110111" => color_data <= "111110110100";
      when "01010111000" => color_data <= "111110110100";
      when "01010111001" => color_data <= "111110110100";
      when "01010111010" => color_data <= "111110110100";
      when "01010111011" => color_data <= "111110110100";
      when "01010111100" => color_data <= "111110110100";
      when "01010111101" => color_data <= "111110110100";
      when "01010111110" => color_data <= "111110110100";
      when "01010111111" => color_data <= "111110110100";
      when "01011000000" => color_data <= "111110110100";
      when "01011000001" => color_data <= "111110110100";
      when "01011000010" => color_data <= "111110110100";
      when "01011000011" => color_data <= "111110110100";
      when "01011000100" => color_data <= "111110110100";
      when "01011000101" => color_data <= "111110110100";
      when "01011000110" => color_data <= "111110110100";
      when "01011000111" => color_data <= "111110110100";
      when "01011001000" => color_data <= "111110110100";
      when "01011001001" => color_data <= "111110110100";
      when "01011001010" => color_data <= "111110110100";
      when "01011001011" => color_data <= "111110110100";
      when "01011001100" => color_data <= "111110110100";
      when "01011001101" => color_data <= "111110110100";
      when "01011001110" => color_data <= "111111010100";
      when "01011001111" => color_data <= "110110100100";
      when "01100000000" => color_data <= "110010100101";
      when "01100000001" => color_data <= "111111100111";
      when "01100000010" => color_data <= "111111010111";
      when "01100000011" => color_data <= "111111010110";
      when "01100000100" => color_data <= "111111010100";
      when "01100000101" => color_data <= "011101100011";
      when "01100000110" => color_data <= "000000010011";
      when "01100000111" => color_data <= "001000110011";
      when "01100001000" => color_data <= "001000110011";
      when "01100001001" => color_data <= "001000110011";
      when "01100001010" => color_data <= "001000110011";
      when "01100001011" => color_data <= "001100110011";
      when "01100001100" => color_data <= "001000110011";
      when "01100001101" => color_data <= "001000110011";
      when "01100001110" => color_data <= "001100110011";
      when "01100001111" => color_data <= "001000110011";
      when "01100010000" => color_data <= "001000110011";
      when "01100010001" => color_data <= "001000110011";
      when "01100010010" => color_data <= "001000110011";
      when "01100010011" => color_data <= "001000110011";
      when "01100010100" => color_data <= "001000110011";
      when "01100010101" => color_data <= "001100110011";
      when "01100010110" => color_data <= "001000110011";
      when "01100010111" => color_data <= "001000110011";
      when "01100011000" => color_data <= "001000110011";
      when "01100011001" => color_data <= "000000100011";
      when "01100011010" => color_data <= "011001010011";
      when "01100011011" => color_data <= "111111010100";
      when "01100011100" => color_data <= "111111000100";
      when "01100011101" => color_data <= "111111000100";
      when "01100011110" => color_data <= "111111000100";
      when "01100011111" => color_data <= "111110110011";
      when "01100100000" => color_data <= "111110110011";
      when "01100100001" => color_data <= "111010110011";
      when "01100100010" => color_data <= "111010110011";
      when "01100100011" => color_data <= "111010110011";
      when "01100100100" => color_data <= "111010110100";
      when "01100100101" => color_data <= "111110110100";
      when "01100100110" => color_data <= "111110110100";
      when "01100100111" => color_data <= "111110110100";
      when "01100101000" => color_data <= "111110110100";
      when "01100101001" => color_data <= "111110110100";
      when "01100101010" => color_data <= "111110110100";
      when "01100101011" => color_data <= "111111000100";
      when "01100101100" => color_data <= "111111000100";
      when "01100101101" => color_data <= "111111000100";
      when "01100101110" => color_data <= "111111000100";
      when "01100101111" => color_data <= "111111000100";
      when "01100110000" => color_data <= "111111000100";
      when "01100110001" => color_data <= "111111000100";
      when "01100110010" => color_data <= "111111000100";
      when "01100110011" => color_data <= "111111000100";
      when "01100110100" => color_data <= "111111000100";
      when "01100110101" => color_data <= "111111000100";
      when "01100110110" => color_data <= "111111000100";
      when "01100110111" => color_data <= "111111000100";
      when "01100111000" => color_data <= "111111000100";
      when "01100111001" => color_data <= "111111000100";
      when "01100111010" => color_data <= "111111000100";
      when "01100111011" => color_data <= "111111000100";
      when "01100111100" => color_data <= "111111000100";
      when "01100111101" => color_data <= "111111000100";
      when "01100111110" => color_data <= "111111000100";
      when "01100111111" => color_data <= "111111000100";
      when "01101000000" => color_data <= "111111000100";
      when "01101000001" => color_data <= "111111000100";
      when "01101000010" => color_data <= "111111000100";
      when "01101000011" => color_data <= "111111000100";
      when "01101000100" => color_data <= "111111000100";
      when "01101000101" => color_data <= "111111000100";
      when "01101000110" => color_data <= "111111000100";
      when "01101000111" => color_data <= "111111000100";
      when "01101001000" => color_data <= "111111000100";
      when "01101001001" => color_data <= "111111000100";
      when "01101001010" => color_data <= "111111000100";
      when "01101001011" => color_data <= "111111000100";
      when "01101001100" => color_data <= "111111000100";
      when "01101001101" => color_data <= "111111000100";
      when "01101001110" => color_data <= "111111010100";
      when "01101001111" => color_data <= "110110100100";
      when "01110000000" => color_data <= "010000110010";
      when "01110000001" => color_data <= "111111100111";
      when "01110000010" => color_data <= "111011000110";
      when "01110000011" => color_data <= "010101000010";
      when "01110000100" => color_data <= "010101000001";
      when "01110000101" => color_data <= "001000100001";
      when "01110000110" => color_data <= "000000000001";
      when "01110000111" => color_data <= "000100010001";
      when "01110001000" => color_data <= "000100010001";
      when "01110001001" => color_data <= "000100010001";
      when "01110001010" => color_data <= "000100010001";
      when "01110001011" => color_data <= "000100010001";
      when "01110001100" => color_data <= "000100010001";
      when "01110001101" => color_data <= "000100010001";
      when "01110001110" => color_data <= "000100010001";
      when "01110001111" => color_data <= "000100010001";
      when "01110010000" => color_data <= "000100010001";
      when "01110010001" => color_data <= "000100010001";
      when "01110010010" => color_data <= "000100010001";
      when "01110010011" => color_data <= "000100010001";
      when "01110010100" => color_data <= "000100010001";
      when "01110010101" => color_data <= "000100010001";
      when "01110010110" => color_data <= "000100010001";
      when "01110010111" => color_data <= "000100010001";
      when "01110011000" => color_data <= "000100010001";
      when "01110011001" => color_data <= "000000000001";
      when "01110011010" => color_data <= "001000100001";
      when "01110011011" => color_data <= "011101010010";
      when "01110011100" => color_data <= "100001100010";
      when "01110011101" => color_data <= "100101110010";
      when "01110011110" => color_data <= "101110000011";
      when "01110011111" => color_data <= "110010010011";
      when "01110100000" => color_data <= "111010100100";
      when "01110100001" => color_data <= "111111000100";
      when "01110100010" => color_data <= "111111000100";
      when "01110100011" => color_data <= "111111000100";
      when "01110100100" => color_data <= "111111000100";
      when "01110100101" => color_data <= "111111000100";
      when "01110100110" => color_data <= "111111000100";
      when "01110100111" => color_data <= "111110110011";
      when "01110101000" => color_data <= "111010110011";
      when "01110101001" => color_data <= "111010110011";
      when "01110101010" => color_data <= "111010110011";
      when "01110101011" => color_data <= "111010110011";
      when "01110101100" => color_data <= "111010110100";
      when "01110101101" => color_data <= "111010110100";
      when "01110101110" => color_data <= "111010110100";
      when "01110101111" => color_data <= "111010110100";
      when "01110110000" => color_data <= "111010110100";
      when "01110110001" => color_data <= "111010110100";
      when "01110110010" => color_data <= "111010110100";
      when "01110110011" => color_data <= "111010110100";
      when "01110110100" => color_data <= "111010110100";
      when "01110110101" => color_data <= "111010110100";
      when "01110110110" => color_data <= "111010110100";
      when "01110110111" => color_data <= "111010110100";
      when "01110111000" => color_data <= "111010110100";
      when "01110111001" => color_data <= "111010110100";
      when "01110111010" => color_data <= "111110110100";
      when "01110111011" => color_data <= "111110110100";
      when "01110111100" => color_data <= "111110110100";
      when "01110111101" => color_data <= "111110110100";
      when "01110111110" => color_data <= "111110110100";
      when "01110111111" => color_data <= "111110110100";
      when "01111000000" => color_data <= "111110110100";
      when "01111000001" => color_data <= "111110110100";
      when "01111000010" => color_data <= "111110110100";
      when "01111000011" => color_data <= "111110110100";
      when "01111000100" => color_data <= "111110110100";
      when "01111000101" => color_data <= "111110110100";
      when "01111000110" => color_data <= "111110110100";
      when "01111000111" => color_data <= "111110110100";
      when "01111001000" => color_data <= "111110110100";
      when "01111001001" => color_data <= "111110110100";
      when "01111001010" => color_data <= "111110110100";
      when "01111001011" => color_data <= "111110110100";
      when "01111001100" => color_data <= "111110110100";
      when "01111001101" => color_data <= "111110110100";
      when "01111001110" => color_data <= "111111010100";
      when "01111001111" => color_data <= "110010010011";
      when "10000000000" => color_data <= "000000000000";
      when "10000000001" => color_data <= "001000100001";
      when "10000000010" => color_data <= "001000010001";
      when "10000000011" => color_data <= "000000000000";
      when "10000000100" => color_data <= "000000000000";
      when "10000000101" => color_data <= "000000000000";
      when "10000000110" => color_data <= "000000000000";
      when "10000000111" => color_data <= "000000000000";
      when "10000001000" => color_data <= "000000000000";
      when "10000001001" => color_data <= "000000000000";
      when "10000001010" => color_data <= "000000000000";
      when "10000001011" => color_data <= "000000000000";
      when "10000001100" => color_data <= "000000000000";
      when "10000001101" => color_data <= "000000000000";
      when "10000001110" => color_data <= "000000000000";
      when "10000001111" => color_data <= "000000000000";
      when "10000010000" => color_data <= "000000000000";
      when "10000010001" => color_data <= "000000000000";
      when "10000010010" => color_data <= "000000000000";
      when "10000010011" => color_data <= "000000000000";
      when "10000010100" => color_data <= "000000000000";
      when "10000010101" => color_data <= "000000000000";
      when "10000010110" => color_data <= "000000000000";
      when "10000010111" => color_data <= "000000000000";
      when "10000011000" => color_data <= "000000000000";
      when "10000011001" => color_data <= "000000000000";
      when "10000011010" => color_data <= "000000000000";
      when "10000011011" => color_data <= "000000000000";
      when "10000011100" => color_data <= "000000000000";
      when "10000011101" => color_data <= "000000000000";
      when "10000011110" => color_data <= "000000000000";
      when "10000011111" => color_data <= "000000000000";
      when "10000100000" => color_data <= "000100010000";
      when "10000100001" => color_data <= "001100110001";
      when "10000100010" => color_data <= "010101000001";
      when "10000100011" => color_data <= "011101010010";
      when "10000100100" => color_data <= "011101100010";
      when "10000100101" => color_data <= "100101110011";
      when "10000100110" => color_data <= "101110010011";
      when "10000100111" => color_data <= "110010100011";
      when "10000101000" => color_data <= "111010110100";
      when "10000101001" => color_data <= "111111000100";
      when "10000101010" => color_data <= "111111000100";
      when "10000101011" => color_data <= "111111000100";
      when "10000101100" => color_data <= "111111000100";
      when "10000101101" => color_data <= "111111000100";
      when "10000101110" => color_data <= "111111000100";
      when "10000101111" => color_data <= "111111000100";
      when "10000110000" => color_data <= "111111000100";
      when "10000110001" => color_data <= "111111000100";
      when "10000110010" => color_data <= "111111000100";
      when "10000110011" => color_data <= "111110110011";
      when "10000110100" => color_data <= "111110110011";
      when "10000110101" => color_data <= "111110110011";
      when "10000110110" => color_data <= "111110110011";
      when "10000110111" => color_data <= "111010110011";
      when "10000111000" => color_data <= "111010100011";
      when "10000111001" => color_data <= "111010100011";
      when "10000111010" => color_data <= "111010100011";
      when "10000111011" => color_data <= "111010100011";
      when "10000111100" => color_data <= "111010100011";
      when "10000111101" => color_data <= "111010100011";
      when "10000111110" => color_data <= "111010100011";
      when "10000111111" => color_data <= "111010100011";
      when "10001000000" => color_data <= "111010100011";
      when "10001000001" => color_data <= "111010100011";
      when "10001000010" => color_data <= "111010100011";
      when "10001000011" => color_data <= "111010100011";
      when "10001000100" => color_data <= "111010100011";
      when "10001000101" => color_data <= "111010100011";
      when "10001000110" => color_data <= "111010100011";
      when "10001000111" => color_data <= "111010100011";
      when "10001001000" => color_data <= "111010100011";
      when "10001001001" => color_data <= "111010100011";
      when "10001001010" => color_data <= "111010100011";
      when "10001001011" => color_data <= "111010100011";
      when "10001001100" => color_data <= "111010100011";
      when "10001001101" => color_data <= "111010100011";
      when "10001001110" => color_data <= "111111010100";
      when "10001001111" => color_data <= "011001010010";
      when "10010000000" => color_data <= "000000000000";
      when "10010000001" => color_data <= "000000000000";
      when "10010000010" => color_data <= "000000000000";
      when "10010000011" => color_data <= "000000000000";
      when "10010000100" => color_data <= "000000000000";
      when "10010000101" => color_data <= "000000000000";
      when "10010000110" => color_data <= "000000000000";
      when "10010000111" => color_data <= "000000000000";
      when "10010001000" => color_data <= "000000000000";
      when "10010001001" => color_data <= "000000000000";
      when "10010001010" => color_data <= "000000000000";
      when "10010001011" => color_data <= "000000000000";
      when "10010001100" => color_data <= "000000000000";
      when "10010001101" => color_data <= "000000000000";
      when "10010001110" => color_data <= "000000000000";
      when "10010001111" => color_data <= "000000000000";
      when "10010010000" => color_data <= "000000000000";
      when "10010010001" => color_data <= "000000000000";
      when "10010010010" => color_data <= "000000000000";
      when "10010010011" => color_data <= "000000000000";
      when "10010010100" => color_data <= "000000000000";
      when "10010010101" => color_data <= "000000000000";
      when "10010010110" => color_data <= "000000000000";
      when "10010010111" => color_data <= "000000000000";
      when "10010011000" => color_data <= "000000000000";
      when "10010011001" => color_data <= "000000000000";
      when "10010011010" => color_data <= "000000000000";
      when "10010011011" => color_data <= "000000000000";
      when "10010011100" => color_data <= "000000000000";
      when "10010011101" => color_data <= "000000000000";
      when "10010011110" => color_data <= "000000000000";
      when "10010011111" => color_data <= "000000000000";
      when "10010100000" => color_data <= "000000000000";
      when "10010100001" => color_data <= "000000000000";
      when "10010100010" => color_data <= "000000000000";
      when "10010100011" => color_data <= "000000000000";
      when "10010100100" => color_data <= "000000000000";
      when "10010100101" => color_data <= "000000000000";
      when "10010100110" => color_data <= "000000000000";
      when "10010100111" => color_data <= "000000000000";
      when "10010101000" => color_data <= "000100010000";
      when "10010101001" => color_data <= "001100110001";
      when "10010101010" => color_data <= "010101000010";
      when "10010101011" => color_data <= "011001010001";
      when "10010101100" => color_data <= "100001100010";
      when "10010101101" => color_data <= "100101100010";
      when "10010101110" => color_data <= "100101110010";
      when "10010101111" => color_data <= "100101110011";
      when "10010110000" => color_data <= "101010000011";
      when "10010110001" => color_data <= "101010000011";
      when "10010110010" => color_data <= "101010000010";
      when "10010110011" => color_data <= "101110000011";
      when "10010110100" => color_data <= "101110010011";
      when "10010110101" => color_data <= "110010010011";
      when "10010110110" => color_data <= "110010010011";
      when "10010110111" => color_data <= "110010010011";
      when "10010111000" => color_data <= "110110100100";
      when "10010111001" => color_data <= "110110100100";
      when "10010111010" => color_data <= "111010110100";
      when "10010111011" => color_data <= "111010100011";
      when "10010111100" => color_data <= "111010100011";
      when "10010111101" => color_data <= "111010100011";
      when "10010111110" => color_data <= "111010100011";
      when "10010111111" => color_data <= "111010100011";
      when "10011000000" => color_data <= "111010100011";
      when "10011000001" => color_data <= "111010100011";
      when "10011000010" => color_data <= "111010100011";
      when "10011000011" => color_data <= "111010100011";
      when "10011000100" => color_data <= "111010100011";
      when "10011000101" => color_data <= "111010100011";
      when "10011000110" => color_data <= "111010100011";
      when "10011000111" => color_data <= "111010100011";
      when "10011001000" => color_data <= "111010100011";
      when "10011001001" => color_data <= "111010100011";
      when "10011001010" => color_data <= "111010100011";
      when "10011001011" => color_data <= "111010100011";
      when "10011001100" => color_data <= "111010110011";
      when "10011001101" => color_data <= "111110110100";
      when "10011001110" => color_data <= "100101110010";
      when "10011001111" => color_data <= "000000000000";
      when others => color_data <= (others => '0');
    end case;
  end process;
end Behavioral;
